module LutMembershipFunctionOnline(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [9:0] i; // @[lut_mem_online.scala 215:18]
  reg  buffer_0; // @[lut_mem_online.scala 219:19]
  reg  buffer_1; // @[lut_mem_online.scala 219:19]
  reg  buffer_2; // @[lut_mem_online.scala 219:19]
  reg  buffer_3; // @[lut_mem_online.scala 219:19]
  reg  buffer_4; // @[lut_mem_online.scala 219:19]
  reg  buffer_5; // @[lut_mem_online.scala 219:19]
  reg  buffer_6; // @[lut_mem_online.scala 219:19]
  reg [4:0] counter; // @[lut_mem_online.scala 221:24]
  reg  outResult; // @[lut_mem_online.scala 224:26]
  wire  _T_2 = counter < 5'ha; // @[lut_mem_online.scala 241:22]
  wire  _GEN_0 = io_inputBit ? 1'h0 : buffer_0; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_1 = i == 10'h0 ? _GEN_0 : buffer_0; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_2 = io_inputBit ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_3 = i == 10'h1 ? _GEN_2 : _GEN_1; // @[lut_mem_online.scala 247:34]
  wire  _GEN_4 = io_inputBit ? 1'h0 : _GEN_3; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_5 = i == 10'h3 ? _GEN_4 : _GEN_3; // @[lut_mem_online.scala 247:34]
  wire  _T_10 = ~io_inputBit; // @[lut_mem_online.scala 249:32]
  wire  _GEN_6 = ~io_inputBit | _GEN_5; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_7 = i == 10'h7 ? _GEN_6 : _GEN_5; // @[lut_mem_online.scala 247:34]
  wire  _GEN_8 = io_inputBit ? 1'h0 : _GEN_7; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_9 = i == 10'h10 ? _GEN_8 : _GEN_7; // @[lut_mem_online.scala 247:34]
  wire  _GEN_10 = ~io_inputBit | _GEN_9; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_11 = i == 10'h21 ? _GEN_10 : _GEN_9; // @[lut_mem_online.scala 247:34]
  wire  _GEN_12 = io_inputBit ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_13 = i == 10'h44 ? _GEN_12 : _GEN_11; // @[lut_mem_online.scala 247:34]
  wire  _GEN_14 = ~io_inputBit | _GEN_13; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_15 = i == 10'h89 ? _GEN_14 : _GEN_13; // @[lut_mem_online.scala 247:34]
  wire  _GEN_16 = ~io_inputBit | _GEN_15; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_17 = i == 10'h114 ? _GEN_16 : _GEN_15; // @[lut_mem_online.scala 247:34]
  wire  _GEN_18 = ~io_inputBit | _GEN_17; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_19 = i == 10'h22a ? _GEN_18 : _GEN_17; // @[lut_mem_online.scala 247:34]
  wire  _GEN_22 = io_inputBit ? 1'h0 : buffer_1; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_23 = i == 10'h0 ? _GEN_22 : buffer_1; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_24 = io_inputBit ? 1'h0 : _GEN_23; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_25 = i == 10'h1 ? _GEN_24 : _GEN_23; // @[lut_mem_online.scala 247:34]
  wire  _GEN_26 = io_inputBit ? 1'h0 : _GEN_25; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_27 = i == 10'h3 ? _GEN_26 : _GEN_25; // @[lut_mem_online.scala 247:34]
  wire  _GEN_28 = ~io_inputBit | _GEN_27; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_29 = i == 10'hf ? _GEN_28 : _GEN_27; // @[lut_mem_online.scala 247:34]
  wire  _GEN_30 = ~io_inputBit | _GEN_29; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_31 = i == 10'h20 ? _GEN_30 : _GEN_29; // @[lut_mem_online.scala 247:34]
  wire  _GEN_32 = ~io_inputBit ? 1'h0 : _GEN_31; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_33 = i == 10'h21 ? _GEN_32 : _GEN_31; // @[lut_mem_online.scala 247:34]
  wire  _GEN_34 = ~io_inputBit | _GEN_33; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_35 = i == 10'h22 ? _GEN_34 : _GEN_33; // @[lut_mem_online.scala 247:34]
  wire  _GEN_36 = io_inputBit ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_37 = i == 10'h42 ? _GEN_36 : _GEN_35; // @[lut_mem_online.scala 247:34]
  wire  _GEN_38 = io_inputBit | _GEN_37; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_39 = i == 10'h44 ? _GEN_38 : _GEN_37; // @[lut_mem_online.scala 247:34]
  wire  _GEN_40 = io_inputBit ? 1'h0 : _GEN_39; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_41 = i == 10'h46 ? _GEN_40 : _GEN_39; // @[lut_mem_online.scala 247:34]
  wire  _GEN_42 = ~io_inputBit | _GEN_41; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_43 = i == 10'h85 ? _GEN_42 : _GEN_41; // @[lut_mem_online.scala 247:34]
  wire  _GEN_44 = ~io_inputBit ? 1'h0 : _GEN_43; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_45 = i == 10'h89 ? _GEN_44 : _GEN_43; // @[lut_mem_online.scala 247:34]
  wire  _GEN_46 = ~io_inputBit | _GEN_45; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_47 = i == 10'h8d ? _GEN_46 : _GEN_45; // @[lut_mem_online.scala 247:34]
  wire  _GEN_48 = ~io_inputBit | _GEN_47; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_49 = i == 10'h10c ? _GEN_48 : _GEN_47; // @[lut_mem_online.scala 247:34]
  wire  _GEN_50 = ~io_inputBit ? 1'h0 : _GEN_49; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_51 = i == 10'h114 ? _GEN_50 : _GEN_49; // @[lut_mem_online.scala 247:34]
  wire  _GEN_52 = ~io_inputBit | _GEN_51; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_53 = i == 10'h11c ? _GEN_52 : _GEN_51; // @[lut_mem_online.scala 247:34]
  wire  _GEN_54 = ~io_inputBit | _GEN_53; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_55 = i == 10'h21a ? _GEN_54 : _GEN_53; // @[lut_mem_online.scala 247:34]
  wire  _GEN_56 = io_inputBit ? 1'h0 : _GEN_55; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_57 = i == 10'h21a ? _GEN_56 : _GEN_55; // @[lut_mem_online.scala 247:34]
  wire  _GEN_58 = ~io_inputBit ? 1'h0 : _GEN_57; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_59 = i == 10'h22a ? _GEN_58 : _GEN_57; // @[lut_mem_online.scala 247:34]
  wire  _GEN_60 = io_inputBit | _GEN_59; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_61 = i == 10'h22a ? _GEN_60 : _GEN_59; // @[lut_mem_online.scala 247:34]
  wire  _GEN_62 = ~io_inputBit | _GEN_61; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_63 = i == 10'h23a ? _GEN_62 : _GEN_61; // @[lut_mem_online.scala 247:34]
  wire  _GEN_66 = io_inputBit ? 1'h0 : buffer_2; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_67 = i == 10'h0 ? _GEN_66 : buffer_2; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_68 = io_inputBit ? 1'h0 : _GEN_67; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_69 = i == 10'h1 ? _GEN_68 : _GEN_67; // @[lut_mem_online.scala 247:34]
  wire  _GEN_70 = io_inputBit ? 1'h0 : _GEN_69; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_71 = i == 10'h8 ? _GEN_70 : _GEN_69; // @[lut_mem_online.scala 247:34]
  wire  _GEN_72 = ~io_inputBit ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_73 = i == 10'hf ? _GEN_72 : _GEN_71; // @[lut_mem_online.scala 247:34]
  wire  _GEN_74 = io_inputBit ? 1'h0 : _GEN_73; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_75 = i == 10'h11 ? _GEN_74 : _GEN_73; // @[lut_mem_online.scala 247:34]
  wire  _GEN_76 = ~io_inputBit ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_77 = i == 10'h20 ? _GEN_76 : _GEN_75; // @[lut_mem_online.scala 247:34]
  wire  _GEN_78 = io_inputBit ? 1'h0 : _GEN_77; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_79 = i == 10'h23 ? _GEN_78 : _GEN_77; // @[lut_mem_online.scala 247:34]
  wire  _GEN_80 = io_inputBit | _GEN_79; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_81 = i == 10'h42 ? _GEN_80 : _GEN_79; // @[lut_mem_online.scala 247:34]
  wire  _GEN_82 = io_inputBit ? 1'h0 : _GEN_81; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_83 = i == 10'h43 ? _GEN_82 : _GEN_81; // @[lut_mem_online.scala 247:34]
  wire  _GEN_84 = io_inputBit | _GEN_83; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_85 = i == 10'h44 ? _GEN_84 : _GEN_83; // @[lut_mem_online.scala 247:34]
  wire  _GEN_86 = io_inputBit ? 1'h0 : _GEN_85; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_87 = i == 10'h45 ? _GEN_86 : _GEN_85; // @[lut_mem_online.scala 247:34]
  wire  _GEN_88 = io_inputBit | _GEN_87; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_89 = i == 10'h46 ? _GEN_88 : _GEN_87; // @[lut_mem_online.scala 247:34]
  wire  _GEN_90 = io_inputBit ? 1'h0 : _GEN_89; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_91 = i == 10'h47 ? _GEN_90 : _GEN_89; // @[lut_mem_online.scala 247:34]
  wire  _GEN_92 = ~io_inputBit ? 1'h0 : _GEN_91; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_93 = i == 10'h85 ? _GEN_92 : _GEN_91; // @[lut_mem_online.scala 247:34]
  wire  _GEN_94 = ~io_inputBit | _GEN_93; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_95 = i == 10'h87 ? _GEN_94 : _GEN_93; // @[lut_mem_online.scala 247:34]
  wire  _GEN_96 = ~io_inputBit ? 1'h0 : _GEN_95; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_97 = i == 10'h89 ? _GEN_96 : _GEN_95; // @[lut_mem_online.scala 247:34]
  wire  _GEN_98 = ~io_inputBit | _GEN_97; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_99 = i == 10'h8b ? _GEN_98 : _GEN_97; // @[lut_mem_online.scala 247:34]
  wire  _GEN_100 = ~io_inputBit ? 1'h0 : _GEN_99; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_101 = i == 10'h8d ? _GEN_100 : _GEN_99; // @[lut_mem_online.scala 247:34]
  wire  _GEN_102 = ~io_inputBit | _GEN_101; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_103 = i == 10'h8f ? _GEN_102 : _GEN_101; // @[lut_mem_online.scala 247:34]
  wire  _GEN_104 = ~io_inputBit ? 1'h0 : _GEN_103; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_105 = i == 10'h10c ? _GEN_104 : _GEN_103; // @[lut_mem_online.scala 247:34]
  wire  _GEN_106 = ~io_inputBit | _GEN_105; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_107 = i == 10'h110 ? _GEN_106 : _GEN_105; // @[lut_mem_online.scala 247:34]
  wire  _GEN_108 = ~io_inputBit ? 1'h0 : _GEN_107; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_109 = i == 10'h114 ? _GEN_108 : _GEN_107; // @[lut_mem_online.scala 247:34]
  wire  _GEN_110 = ~io_inputBit | _GEN_109; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_111 = i == 10'h118 ? _GEN_110 : _GEN_109; // @[lut_mem_online.scala 247:34]
  wire  _GEN_112 = ~io_inputBit ? 1'h0 : _GEN_111; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_113 = i == 10'h11c ? _GEN_112 : _GEN_111; // @[lut_mem_online.scala 247:34]
  wire  _GEN_114 = ~io_inputBit | _GEN_113; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_115 = i == 10'h120 ? _GEN_114 : _GEN_113; // @[lut_mem_online.scala 247:34]
  wire  _GEN_116 = ~io_inputBit ? 1'h0 : _GEN_115; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_117 = i == 10'h21a ? _GEN_116 : _GEN_115; // @[lut_mem_online.scala 247:34]
  wire  _GEN_118 = io_inputBit | _GEN_117; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_119 = i == 10'h21a ? _GEN_118 : _GEN_117; // @[lut_mem_online.scala 247:34]
  wire  _GEN_120 = ~io_inputBit | _GEN_119; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_121 = i == 10'h222 ? _GEN_120 : _GEN_119; // @[lut_mem_online.scala 247:34]
  wire  _GEN_122 = io_inputBit ? 1'h0 : _GEN_121; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_123 = i == 10'h222 ? _GEN_122 : _GEN_121; // @[lut_mem_online.scala 247:34]
  wire  _GEN_124 = ~io_inputBit ? 1'h0 : _GEN_123; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_125 = i == 10'h22a ? _GEN_124 : _GEN_123; // @[lut_mem_online.scala 247:34]
  wire  _GEN_126 = io_inputBit | _GEN_125; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_127 = i == 10'h22a ? _GEN_126 : _GEN_125; // @[lut_mem_online.scala 247:34]
  wire  _GEN_128 = ~io_inputBit | _GEN_127; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_129 = i == 10'h232 ? _GEN_128 : _GEN_127; // @[lut_mem_online.scala 247:34]
  wire  _GEN_130 = io_inputBit ? 1'h0 : _GEN_129; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_131 = i == 10'h232 ? _GEN_130 : _GEN_129; // @[lut_mem_online.scala 247:34]
  wire  _GEN_132 = ~io_inputBit ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_133 = i == 10'h23a ? _GEN_132 : _GEN_131; // @[lut_mem_online.scala 247:34]
  wire  _GEN_134 = io_inputBit | _GEN_133; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_135 = i == 10'h23a ? _GEN_134 : _GEN_133; // @[lut_mem_online.scala 247:34]
  wire  _GEN_136 = ~io_inputBit | _GEN_135; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_137 = i == 10'h242 ? _GEN_136 : _GEN_135; // @[lut_mem_online.scala 247:34]
  wire  _GEN_140 = io_inputBit ? 1'h0 : buffer_3; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_141 = i == 10'h0 ? _GEN_140 : buffer_3; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_142 = io_inputBit ? 1'h0 : _GEN_141; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_143 = i == 10'h1 ? _GEN_142 : _GEN_141; // @[lut_mem_online.scala 247:34]
  wire  _GEN_144 = io_inputBit ? 1'h0 : _GEN_143; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_145 = i == 10'h8 ? _GEN_144 : _GEN_143; // @[lut_mem_online.scala 247:34]
  wire  _GEN_146 = ~io_inputBit ? 1'h0 : _GEN_145; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_147 = i == 10'hf ? _GEN_146 : _GEN_145; // @[lut_mem_online.scala 247:34]
  wire  _GEN_148 = io_inputBit ? 1'h0 : _GEN_147; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_149 = i == 10'h11 ? _GEN_148 : _GEN_147; // @[lut_mem_online.scala 247:34]
  wire  _GEN_150 = ~io_inputBit ? 1'h0 : _GEN_149; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_151 = i == 10'h20 ? _GEN_150 : _GEN_149; // @[lut_mem_online.scala 247:34]
  wire  _GEN_152 = io_inputBit ? 1'h0 : _GEN_151; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_153 = i == 10'h23 ? _GEN_152 : _GEN_151; // @[lut_mem_online.scala 247:34]
  wire  _GEN_154 = ~io_inputBit ? 1'h0 : _GEN_153; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_155 = i == 10'h85 ? _GEN_154 : _GEN_153; // @[lut_mem_online.scala 247:34]
  wire  _GEN_156 = ~io_inputBit | _GEN_155; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_157 = i == 10'h86 ? _GEN_156 : _GEN_155; // @[lut_mem_online.scala 247:34]
  wire  _GEN_158 = ~io_inputBit ? 1'h0 : _GEN_157; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_159 = i == 10'h87 ? _GEN_158 : _GEN_157; // @[lut_mem_online.scala 247:34]
  wire  _GEN_160 = ~io_inputBit | _GEN_159; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_161 = i == 10'h88 ? _GEN_160 : _GEN_159; // @[lut_mem_online.scala 247:34]
  wire  _GEN_162 = ~io_inputBit ? 1'h0 : _GEN_161; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_163 = i == 10'h89 ? _GEN_162 : _GEN_161; // @[lut_mem_online.scala 247:34]
  wire  _GEN_164 = ~io_inputBit | _GEN_163; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_165 = i == 10'h8a ? _GEN_164 : _GEN_163; // @[lut_mem_online.scala 247:34]
  wire  _GEN_166 = ~io_inputBit ? 1'h0 : _GEN_165; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_167 = i == 10'h8b ? _GEN_166 : _GEN_165; // @[lut_mem_online.scala 247:34]
  wire  _GEN_168 = ~io_inputBit | _GEN_167; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_169 = i == 10'h8c ? _GEN_168 : _GEN_167; // @[lut_mem_online.scala 247:34]
  wire  _GEN_170 = ~io_inputBit ? 1'h0 : _GEN_169; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_171 = i == 10'h8d ? _GEN_170 : _GEN_169; // @[lut_mem_online.scala 247:34]
  wire  _GEN_172 = ~io_inputBit | _GEN_171; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_173 = i == 10'h8e ? _GEN_172 : _GEN_171; // @[lut_mem_online.scala 247:34]
  wire  _GEN_174 = ~io_inputBit ? 1'h0 : _GEN_173; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_175 = i == 10'h8f ? _GEN_174 : _GEN_173; // @[lut_mem_online.scala 247:34]
  wire  _GEN_176 = ~io_inputBit | _GEN_175; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_177 = i == 10'h90 ? _GEN_176 : _GEN_175; // @[lut_mem_online.scala 247:34]
  wire  _GEN_178 = ~io_inputBit ? 1'h0 : _GEN_177; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_179 = i == 10'h10c ? _GEN_178 : _GEN_177; // @[lut_mem_online.scala 247:34]
  wire  _GEN_180 = ~io_inputBit | _GEN_179; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_181 = i == 10'h10e ? _GEN_180 : _GEN_179; // @[lut_mem_online.scala 247:34]
  wire  _GEN_182 = ~io_inputBit ? 1'h0 : _GEN_181; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_183 = i == 10'h110 ? _GEN_182 : _GEN_181; // @[lut_mem_online.scala 247:34]
  wire  _GEN_184 = ~io_inputBit | _GEN_183; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_185 = i == 10'h112 ? _GEN_184 : _GEN_183; // @[lut_mem_online.scala 247:34]
  wire  _GEN_186 = ~io_inputBit ? 1'h0 : _GEN_185; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_187 = i == 10'h114 ? _GEN_186 : _GEN_185; // @[lut_mem_online.scala 247:34]
  wire  _GEN_188 = ~io_inputBit | _GEN_187; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_189 = i == 10'h116 ? _GEN_188 : _GEN_187; // @[lut_mem_online.scala 247:34]
  wire  _GEN_190 = ~io_inputBit ? 1'h0 : _GEN_189; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_191 = i == 10'h118 ? _GEN_190 : _GEN_189; // @[lut_mem_online.scala 247:34]
  wire  _GEN_192 = ~io_inputBit | _GEN_191; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_193 = i == 10'h11a ? _GEN_192 : _GEN_191; // @[lut_mem_online.scala 247:34]
  wire  _GEN_194 = ~io_inputBit ? 1'h0 : _GEN_193; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_195 = i == 10'h11c ? _GEN_194 : _GEN_193; // @[lut_mem_online.scala 247:34]
  wire  _GEN_196 = ~io_inputBit | _GEN_195; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_197 = i == 10'h11e ? _GEN_196 : _GEN_195; // @[lut_mem_online.scala 247:34]
  wire  _GEN_198 = ~io_inputBit ? 1'h0 : _GEN_197; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_199 = i == 10'h120 ? _GEN_198 : _GEN_197; // @[lut_mem_online.scala 247:34]
  wire  _GEN_200 = ~io_inputBit | _GEN_199; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_201 = i == 10'h122 ? _GEN_200 : _GEN_199; // @[lut_mem_online.scala 247:34]
  wire  _GEN_202 = ~io_inputBit ? 1'h0 : _GEN_201; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_203 = i == 10'h21a ? _GEN_202 : _GEN_201; // @[lut_mem_online.scala 247:34]
  wire  _GEN_204 = io_inputBit | _GEN_203; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_205 = i == 10'h21a ? _GEN_204 : _GEN_203; // @[lut_mem_online.scala 247:34]
  wire  _GEN_206 = ~io_inputBit | _GEN_205; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_207 = i == 10'h21e ? _GEN_206 : _GEN_205; // @[lut_mem_online.scala 247:34]
  wire  _GEN_208 = io_inputBit ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_209 = i == 10'h21e ? _GEN_208 : _GEN_207; // @[lut_mem_online.scala 247:34]
  wire  _GEN_210 = ~io_inputBit ? 1'h0 : _GEN_209; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_211 = i == 10'h222 ? _GEN_210 : _GEN_209; // @[lut_mem_online.scala 247:34]
  wire  _GEN_212 = io_inputBit | _GEN_211; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_213 = i == 10'h222 ? _GEN_212 : _GEN_211; // @[lut_mem_online.scala 247:34]
  wire  _GEN_214 = ~io_inputBit | _GEN_213; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_215 = i == 10'h226 ? _GEN_214 : _GEN_213; // @[lut_mem_online.scala 247:34]
  wire  _GEN_216 = io_inputBit ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_217 = i == 10'h226 ? _GEN_216 : _GEN_215; // @[lut_mem_online.scala 247:34]
  wire  _GEN_218 = ~io_inputBit ? 1'h0 : _GEN_217; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_219 = i == 10'h22a ? _GEN_218 : _GEN_217; // @[lut_mem_online.scala 247:34]
  wire  _GEN_220 = io_inputBit | _GEN_219; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_221 = i == 10'h22a ? _GEN_220 : _GEN_219; // @[lut_mem_online.scala 247:34]
  wire  _GEN_222 = ~io_inputBit | _GEN_221; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_223 = i == 10'h22e ? _GEN_222 : _GEN_221; // @[lut_mem_online.scala 247:34]
  wire  _GEN_224 = io_inputBit ? 1'h0 : _GEN_223; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_225 = i == 10'h22e ? _GEN_224 : _GEN_223; // @[lut_mem_online.scala 247:34]
  wire  _GEN_226 = ~io_inputBit ? 1'h0 : _GEN_225; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_227 = i == 10'h232 ? _GEN_226 : _GEN_225; // @[lut_mem_online.scala 247:34]
  wire  _GEN_228 = io_inputBit | _GEN_227; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_229 = i == 10'h232 ? _GEN_228 : _GEN_227; // @[lut_mem_online.scala 247:34]
  wire  _GEN_230 = ~io_inputBit | _GEN_229; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_231 = i == 10'h236 ? _GEN_230 : _GEN_229; // @[lut_mem_online.scala 247:34]
  wire  _GEN_232 = io_inputBit ? 1'h0 : _GEN_231; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_233 = i == 10'h236 ? _GEN_232 : _GEN_231; // @[lut_mem_online.scala 247:34]
  wire  _GEN_234 = ~io_inputBit ? 1'h0 : _GEN_233; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_235 = i == 10'h23a ? _GEN_234 : _GEN_233; // @[lut_mem_online.scala 247:34]
  wire  _GEN_236 = io_inputBit | _GEN_235; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_237 = i == 10'h23a ? _GEN_236 : _GEN_235; // @[lut_mem_online.scala 247:34]
  wire  _GEN_238 = ~io_inputBit | _GEN_237; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_239 = i == 10'h23e ? _GEN_238 : _GEN_237; // @[lut_mem_online.scala 247:34]
  wire  _GEN_240 = io_inputBit ? 1'h0 : _GEN_239; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_241 = i == 10'h23e ? _GEN_240 : _GEN_239; // @[lut_mem_online.scala 247:34]
  wire  _GEN_242 = ~io_inputBit ? 1'h0 : _GEN_241; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_243 = i == 10'h242 ? _GEN_242 : _GEN_241; // @[lut_mem_online.scala 247:34]
  wire  _GEN_244 = io_inputBit | _GEN_243; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_245 = i == 10'h242 ? _GEN_244 : _GEN_243; // @[lut_mem_online.scala 247:34]
  wire  _GEN_246 = ~io_inputBit | _GEN_245; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_247 = i == 10'h246 ? _GEN_246 : _GEN_245; // @[lut_mem_online.scala 247:34]
  wire  _GEN_250 = io_inputBit ? 1'h0 : buffer_4; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_251 = i == 10'h0 ? _GEN_250 : buffer_4; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_252 = io_inputBit ? 1'h0 : _GEN_251; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_253 = i == 10'h1 ? _GEN_252 : _GEN_251; // @[lut_mem_online.scala 247:34]
  wire  _GEN_254 = io_inputBit ? 1'h0 : _GEN_253; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_255 = i == 10'h8 ? _GEN_254 : _GEN_253; // @[lut_mem_online.scala 247:34]
  wire  _GEN_256 = ~io_inputBit | _GEN_255; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_257 = i == 10'hf ? _GEN_256 : _GEN_255; // @[lut_mem_online.scala 247:34]
  wire  _GEN_258 = io_inputBit ? 1'h0 : _GEN_257; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_259 = i == 10'h11 ? _GEN_258 : _GEN_257; // @[lut_mem_online.scala 247:34]
  wire  _GEN_260 = ~io_inputBit | _GEN_259; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_261 = i == 10'h20 ? _GEN_260 : _GEN_259; // @[lut_mem_online.scala 247:34]
  wire  _GEN_262 = io_inputBit ? 1'h0 : _GEN_261; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_263 = i == 10'h48 ? _GEN_262 : _GEN_261; // @[lut_mem_online.scala 247:34]
  wire  _GEN_264 = io_inputBit ? 1'h0 : _GEN_263; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_265 = i == 10'h91 ? _GEN_264 : _GEN_263; // @[lut_mem_online.scala 247:34]
  wire  _GEN_266 = ~io_inputBit | _GEN_265; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_267 = i == 10'h10b ? _GEN_266 : _GEN_265; // @[lut_mem_online.scala 247:34]
  wire  _GEN_268 = ~io_inputBit ? 1'h0 : _GEN_267; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_269 = i == 10'h10c ? _GEN_268 : _GEN_267; // @[lut_mem_online.scala 247:34]
  wire  _GEN_270 = ~io_inputBit | _GEN_269; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_271 = i == 10'h10d ? _GEN_270 : _GEN_269; // @[lut_mem_online.scala 247:34]
  wire  _GEN_272 = ~io_inputBit ? 1'h0 : _GEN_271; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_273 = i == 10'h10e ? _GEN_272 : _GEN_271; // @[lut_mem_online.scala 247:34]
  wire  _GEN_274 = ~io_inputBit | _GEN_273; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_275 = i == 10'h10f ? _GEN_274 : _GEN_273; // @[lut_mem_online.scala 247:34]
  wire  _GEN_276 = ~io_inputBit ? 1'h0 : _GEN_275; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_277 = i == 10'h110 ? _GEN_276 : _GEN_275; // @[lut_mem_online.scala 247:34]
  wire  _GEN_278 = ~io_inputBit | _GEN_277; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_279 = i == 10'h111 ? _GEN_278 : _GEN_277; // @[lut_mem_online.scala 247:34]
  wire  _GEN_280 = ~io_inputBit ? 1'h0 : _GEN_279; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_281 = i == 10'h112 ? _GEN_280 : _GEN_279; // @[lut_mem_online.scala 247:34]
  wire  _GEN_282 = ~io_inputBit | _GEN_281; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_283 = i == 10'h113 ? _GEN_282 : _GEN_281; // @[lut_mem_online.scala 247:34]
  wire  _GEN_284 = ~io_inputBit ? 1'h0 : _GEN_283; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_285 = i == 10'h114 ? _GEN_284 : _GEN_283; // @[lut_mem_online.scala 247:34]
  wire  _GEN_286 = ~io_inputBit | _GEN_285; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_287 = i == 10'h115 ? _GEN_286 : _GEN_285; // @[lut_mem_online.scala 247:34]
  wire  _GEN_288 = ~io_inputBit ? 1'h0 : _GEN_287; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_289 = i == 10'h116 ? _GEN_288 : _GEN_287; // @[lut_mem_online.scala 247:34]
  wire  _GEN_290 = ~io_inputBit | _GEN_289; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_291 = i == 10'h117 ? _GEN_290 : _GEN_289; // @[lut_mem_online.scala 247:34]
  wire  _GEN_292 = ~io_inputBit ? 1'h0 : _GEN_291; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_293 = i == 10'h118 ? _GEN_292 : _GEN_291; // @[lut_mem_online.scala 247:34]
  wire  _GEN_294 = ~io_inputBit | _GEN_293; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_295 = i == 10'h119 ? _GEN_294 : _GEN_293; // @[lut_mem_online.scala 247:34]
  wire  _GEN_296 = ~io_inputBit ? 1'h0 : _GEN_295; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_297 = i == 10'h11a ? _GEN_296 : _GEN_295; // @[lut_mem_online.scala 247:34]
  wire  _GEN_298 = ~io_inputBit | _GEN_297; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_299 = i == 10'h11b ? _GEN_298 : _GEN_297; // @[lut_mem_online.scala 247:34]
  wire  _GEN_300 = ~io_inputBit ? 1'h0 : _GEN_299; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_301 = i == 10'h11c ? _GEN_300 : _GEN_299; // @[lut_mem_online.scala 247:34]
  wire  _GEN_302 = ~io_inputBit | _GEN_301; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_303 = i == 10'h11d ? _GEN_302 : _GEN_301; // @[lut_mem_online.scala 247:34]
  wire  _GEN_304 = ~io_inputBit ? 1'h0 : _GEN_303; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_305 = i == 10'h11e ? _GEN_304 : _GEN_303; // @[lut_mem_online.scala 247:34]
  wire  _GEN_306 = ~io_inputBit | _GEN_305; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_307 = i == 10'h11f ? _GEN_306 : _GEN_305; // @[lut_mem_online.scala 247:34]
  wire  _GEN_308 = ~io_inputBit ? 1'h0 : _GEN_307; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_309 = i == 10'h120 ? _GEN_308 : _GEN_307; // @[lut_mem_online.scala 247:34]
  wire  _GEN_310 = ~io_inputBit | _GEN_309; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_311 = i == 10'h121 ? _GEN_310 : _GEN_309; // @[lut_mem_online.scala 247:34]
  wire  _GEN_312 = ~io_inputBit ? 1'h0 : _GEN_311; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_313 = i == 10'h122 ? _GEN_312 : _GEN_311; // @[lut_mem_online.scala 247:34]
  wire  _GEN_314 = ~io_inputBit | _GEN_313; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_315 = i == 10'h123 ? _GEN_314 : _GEN_313; // @[lut_mem_online.scala 247:34]
  wire  _GEN_316 = ~io_inputBit | _GEN_315; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_317 = i == 10'h218 ? _GEN_316 : _GEN_315; // @[lut_mem_online.scala 247:34]
  wire  _GEN_318 = io_inputBit ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_319 = i == 10'h218 ? _GEN_318 : _GEN_317; // @[lut_mem_online.scala 247:34]
  wire  _GEN_320 = ~io_inputBit ? 1'h0 : _GEN_319; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_321 = i == 10'h21a ? _GEN_320 : _GEN_319; // @[lut_mem_online.scala 247:34]
  wire  _GEN_322 = io_inputBit | _GEN_321; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_323 = i == 10'h21a ? _GEN_322 : _GEN_321; // @[lut_mem_online.scala 247:34]
  wire  _GEN_324 = ~io_inputBit | _GEN_323; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_325 = i == 10'h21c ? _GEN_324 : _GEN_323; // @[lut_mem_online.scala 247:34]
  wire  _GEN_326 = io_inputBit ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_327 = i == 10'h21c ? _GEN_326 : _GEN_325; // @[lut_mem_online.scala 247:34]
  wire  _GEN_328 = ~io_inputBit ? 1'h0 : _GEN_327; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_329 = i == 10'h21e ? _GEN_328 : _GEN_327; // @[lut_mem_online.scala 247:34]
  wire  _GEN_330 = io_inputBit | _GEN_329; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_331 = i == 10'h21e ? _GEN_330 : _GEN_329; // @[lut_mem_online.scala 247:34]
  wire  _GEN_332 = ~io_inputBit | _GEN_331; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_333 = i == 10'h220 ? _GEN_332 : _GEN_331; // @[lut_mem_online.scala 247:34]
  wire  _GEN_334 = io_inputBit ? 1'h0 : _GEN_333; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_335 = i == 10'h220 ? _GEN_334 : _GEN_333; // @[lut_mem_online.scala 247:34]
  wire  _GEN_336 = ~io_inputBit ? 1'h0 : _GEN_335; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_337 = i == 10'h222 ? _GEN_336 : _GEN_335; // @[lut_mem_online.scala 247:34]
  wire  _GEN_338 = io_inputBit | _GEN_337; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_339 = i == 10'h222 ? _GEN_338 : _GEN_337; // @[lut_mem_online.scala 247:34]
  wire  _GEN_340 = ~io_inputBit | _GEN_339; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_341 = i == 10'h224 ? _GEN_340 : _GEN_339; // @[lut_mem_online.scala 247:34]
  wire  _GEN_342 = io_inputBit ? 1'h0 : _GEN_341; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_343 = i == 10'h224 ? _GEN_342 : _GEN_341; // @[lut_mem_online.scala 247:34]
  wire  _GEN_344 = ~io_inputBit ? 1'h0 : _GEN_343; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_345 = i == 10'h226 ? _GEN_344 : _GEN_343; // @[lut_mem_online.scala 247:34]
  wire  _GEN_346 = io_inputBit | _GEN_345; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_347 = i == 10'h226 ? _GEN_346 : _GEN_345; // @[lut_mem_online.scala 247:34]
  wire  _GEN_348 = ~io_inputBit | _GEN_347; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_349 = i == 10'h228 ? _GEN_348 : _GEN_347; // @[lut_mem_online.scala 247:34]
  wire  _GEN_350 = io_inputBit ? 1'h0 : _GEN_349; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_351 = i == 10'h228 ? _GEN_350 : _GEN_349; // @[lut_mem_online.scala 247:34]
  wire  _GEN_352 = ~io_inputBit ? 1'h0 : _GEN_351; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_353 = i == 10'h22a ? _GEN_352 : _GEN_351; // @[lut_mem_online.scala 247:34]
  wire  _GEN_354 = io_inputBit | _GEN_353; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_355 = i == 10'h22a ? _GEN_354 : _GEN_353; // @[lut_mem_online.scala 247:34]
  wire  _GEN_356 = ~io_inputBit | _GEN_355; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_357 = i == 10'h22c ? _GEN_356 : _GEN_355; // @[lut_mem_online.scala 247:34]
  wire  _GEN_358 = io_inputBit ? 1'h0 : _GEN_357; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_359 = i == 10'h22c ? _GEN_358 : _GEN_357; // @[lut_mem_online.scala 247:34]
  wire  _GEN_360 = ~io_inputBit ? 1'h0 : _GEN_359; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_361 = i == 10'h22e ? _GEN_360 : _GEN_359; // @[lut_mem_online.scala 247:34]
  wire  _GEN_362 = io_inputBit | _GEN_361; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_363 = i == 10'h22e ? _GEN_362 : _GEN_361; // @[lut_mem_online.scala 247:34]
  wire  _GEN_364 = ~io_inputBit | _GEN_363; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_365 = i == 10'h230 ? _GEN_364 : _GEN_363; // @[lut_mem_online.scala 247:34]
  wire  _GEN_366 = io_inputBit ? 1'h0 : _GEN_365; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_367 = i == 10'h230 ? _GEN_366 : _GEN_365; // @[lut_mem_online.scala 247:34]
  wire  _GEN_368 = ~io_inputBit ? 1'h0 : _GEN_367; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_369 = i == 10'h232 ? _GEN_368 : _GEN_367; // @[lut_mem_online.scala 247:34]
  wire  _GEN_370 = io_inputBit | _GEN_369; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_371 = i == 10'h232 ? _GEN_370 : _GEN_369; // @[lut_mem_online.scala 247:34]
  wire  _GEN_372 = ~io_inputBit | _GEN_371; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_373 = i == 10'h234 ? _GEN_372 : _GEN_371; // @[lut_mem_online.scala 247:34]
  wire  _GEN_374 = io_inputBit ? 1'h0 : _GEN_373; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_375 = i == 10'h234 ? _GEN_374 : _GEN_373; // @[lut_mem_online.scala 247:34]
  wire  _GEN_376 = ~io_inputBit ? 1'h0 : _GEN_375; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_377 = i == 10'h236 ? _GEN_376 : _GEN_375; // @[lut_mem_online.scala 247:34]
  wire  _GEN_378 = io_inputBit | _GEN_377; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_379 = i == 10'h236 ? _GEN_378 : _GEN_377; // @[lut_mem_online.scala 247:34]
  wire  _GEN_380 = ~io_inputBit | _GEN_379; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_381 = i == 10'h238 ? _GEN_380 : _GEN_379; // @[lut_mem_online.scala 247:34]
  wire  _GEN_382 = io_inputBit ? 1'h0 : _GEN_381; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_383 = i == 10'h238 ? _GEN_382 : _GEN_381; // @[lut_mem_online.scala 247:34]
  wire  _GEN_384 = ~io_inputBit ? 1'h0 : _GEN_383; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_385 = i == 10'h23a ? _GEN_384 : _GEN_383; // @[lut_mem_online.scala 247:34]
  wire  _GEN_386 = io_inputBit | _GEN_385; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_387 = i == 10'h23a ? _GEN_386 : _GEN_385; // @[lut_mem_online.scala 247:34]
  wire  _GEN_388 = ~io_inputBit | _GEN_387; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_389 = i == 10'h23c ? _GEN_388 : _GEN_387; // @[lut_mem_online.scala 247:34]
  wire  _GEN_390 = io_inputBit ? 1'h0 : _GEN_389; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_391 = i == 10'h23c ? _GEN_390 : _GEN_389; // @[lut_mem_online.scala 247:34]
  wire  _GEN_392 = ~io_inputBit ? 1'h0 : _GEN_391; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_393 = i == 10'h23e ? _GEN_392 : _GEN_391; // @[lut_mem_online.scala 247:34]
  wire  _GEN_394 = io_inputBit | _GEN_393; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_395 = i == 10'h23e ? _GEN_394 : _GEN_393; // @[lut_mem_online.scala 247:34]
  wire  _GEN_396 = ~io_inputBit | _GEN_395; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_397 = i == 10'h240 ? _GEN_396 : _GEN_395; // @[lut_mem_online.scala 247:34]
  wire  _GEN_398 = io_inputBit ? 1'h0 : _GEN_397; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_399 = i == 10'h240 ? _GEN_398 : _GEN_397; // @[lut_mem_online.scala 247:34]
  wire  _GEN_400 = ~io_inputBit ? 1'h0 : _GEN_399; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_401 = i == 10'h242 ? _GEN_400 : _GEN_399; // @[lut_mem_online.scala 247:34]
  wire  _GEN_402 = io_inputBit | _GEN_401; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_403 = i == 10'h242 ? _GEN_402 : _GEN_401; // @[lut_mem_online.scala 247:34]
  wire  _GEN_404 = ~io_inputBit | _GEN_403; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_405 = i == 10'h244 ? _GEN_404 : _GEN_403; // @[lut_mem_online.scala 247:34]
  wire  _GEN_406 = io_inputBit ? 1'h0 : _GEN_405; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_407 = i == 10'h244 ? _GEN_406 : _GEN_405; // @[lut_mem_online.scala 247:34]
  wire  _GEN_408 = ~io_inputBit ? 1'h0 : _GEN_407; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_409 = i == 10'h246 ? _GEN_408 : _GEN_407; // @[lut_mem_online.scala 247:34]
  wire  _GEN_410 = io_inputBit | _GEN_409; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_411 = i == 10'h246 ? _GEN_410 : _GEN_409; // @[lut_mem_online.scala 247:34]
  wire  _GEN_412 = ~io_inputBit | _GEN_411; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_413 = i == 10'h248 ? _GEN_412 : _GEN_411; // @[lut_mem_online.scala 247:34]
  wire  _GEN_416 = io_inputBit ? 1'h0 : buffer_5; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_417 = i == 10'h0 ? _GEN_416 : buffer_5; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_418 = io_inputBit ? 1'h0 : _GEN_417; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_419 = i == 10'h1 ? _GEN_418 : _GEN_417; // @[lut_mem_online.scala 247:34]
  wire  _GEN_420 = io_inputBit ? 1'h0 : _GEN_419; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_421 = i == 10'h8 ? _GEN_420 : _GEN_419; // @[lut_mem_online.scala 247:34]
  wire  _GEN_422 = ~io_inputBit ? 1'h0 : _GEN_421; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_423 = i == 10'hf ? _GEN_422 : _GEN_421; // @[lut_mem_online.scala 247:34]
  wire  _GEN_424 = io_inputBit ? 1'h0 : _GEN_423; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_425 = i == 10'h11 ? _GEN_424 : _GEN_423; // @[lut_mem_online.scala 247:34]
  wire  _GEN_426 = ~io_inputBit ? 1'h0 : _GEN_425; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_427 = i == 10'h20 ? _GEN_426 : _GEN_425; // @[lut_mem_online.scala 247:34]
  wire  _GEN_428 = io_inputBit ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_429 = i == 10'h48 ? _GEN_428 : _GEN_427; // @[lut_mem_online.scala 247:34]
  wire  _GEN_430 = ~io_inputBit ? 1'h0 : _GEN_429; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_431 = i == 10'h10b ? _GEN_430 : _GEN_429; // @[lut_mem_online.scala 247:34]
  wire  _GEN_432 = io_inputBit ? 1'h0 : _GEN_431; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_433 = i == 10'h124 ? _GEN_432 : _GEN_431; // @[lut_mem_online.scala 247:34]
  wire  _GEN_434 = ~io_inputBit ? 1'h0 : _GEN_433; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_435 = i == 10'h218 ? _GEN_434 : _GEN_433; // @[lut_mem_online.scala 247:34]
  wire  _GEN_436 = io_inputBit | _GEN_435; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_437 = i == 10'h218 ? _GEN_436 : _GEN_435; // @[lut_mem_online.scala 247:34]
  wire  _GEN_438 = ~io_inputBit | _GEN_437; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_439 = i == 10'h219 ? _GEN_438 : _GEN_437; // @[lut_mem_online.scala 247:34]
  wire  _GEN_440 = io_inputBit ? 1'h0 : _GEN_439; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_441 = i == 10'h219 ? _GEN_440 : _GEN_439; // @[lut_mem_online.scala 247:34]
  wire  _GEN_442 = ~io_inputBit ? 1'h0 : _GEN_441; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_443 = i == 10'h21a ? _GEN_442 : _GEN_441; // @[lut_mem_online.scala 247:34]
  wire  _GEN_444 = io_inputBit | _GEN_443; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_445 = i == 10'h21a ? _GEN_444 : _GEN_443; // @[lut_mem_online.scala 247:34]
  wire  _GEN_446 = ~io_inputBit | _GEN_445; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_447 = i == 10'h21b ? _GEN_446 : _GEN_445; // @[lut_mem_online.scala 247:34]
  wire  _GEN_448 = io_inputBit ? 1'h0 : _GEN_447; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_449 = i == 10'h21b ? _GEN_448 : _GEN_447; // @[lut_mem_online.scala 247:34]
  wire  _GEN_450 = ~io_inputBit ? 1'h0 : _GEN_449; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_451 = i == 10'h21c ? _GEN_450 : _GEN_449; // @[lut_mem_online.scala 247:34]
  wire  _GEN_452 = io_inputBit | _GEN_451; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_453 = i == 10'h21c ? _GEN_452 : _GEN_451; // @[lut_mem_online.scala 247:34]
  wire  _GEN_454 = ~io_inputBit | _GEN_453; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_455 = i == 10'h21d ? _GEN_454 : _GEN_453; // @[lut_mem_online.scala 247:34]
  wire  _GEN_456 = io_inputBit ? 1'h0 : _GEN_455; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_457 = i == 10'h21d ? _GEN_456 : _GEN_455; // @[lut_mem_online.scala 247:34]
  wire  _GEN_458 = ~io_inputBit ? 1'h0 : _GEN_457; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_459 = i == 10'h21e ? _GEN_458 : _GEN_457; // @[lut_mem_online.scala 247:34]
  wire  _GEN_460 = io_inputBit | _GEN_459; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_461 = i == 10'h21e ? _GEN_460 : _GEN_459; // @[lut_mem_online.scala 247:34]
  wire  _GEN_462 = ~io_inputBit | _GEN_461; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_463 = i == 10'h21f ? _GEN_462 : _GEN_461; // @[lut_mem_online.scala 247:34]
  wire  _GEN_464 = io_inputBit ? 1'h0 : _GEN_463; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_465 = i == 10'h21f ? _GEN_464 : _GEN_463; // @[lut_mem_online.scala 247:34]
  wire  _GEN_466 = ~io_inputBit ? 1'h0 : _GEN_465; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_467 = i == 10'h220 ? _GEN_466 : _GEN_465; // @[lut_mem_online.scala 247:34]
  wire  _GEN_468 = io_inputBit | _GEN_467; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_469 = i == 10'h220 ? _GEN_468 : _GEN_467; // @[lut_mem_online.scala 247:34]
  wire  _GEN_470 = ~io_inputBit | _GEN_469; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_471 = i == 10'h221 ? _GEN_470 : _GEN_469; // @[lut_mem_online.scala 247:34]
  wire  _GEN_472 = io_inputBit ? 1'h0 : _GEN_471; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_473 = i == 10'h221 ? _GEN_472 : _GEN_471; // @[lut_mem_online.scala 247:34]
  wire  _GEN_474 = ~io_inputBit ? 1'h0 : _GEN_473; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_475 = i == 10'h222 ? _GEN_474 : _GEN_473; // @[lut_mem_online.scala 247:34]
  wire  _GEN_476 = io_inputBit | _GEN_475; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_477 = i == 10'h222 ? _GEN_476 : _GEN_475; // @[lut_mem_online.scala 247:34]
  wire  _GEN_478 = ~io_inputBit | _GEN_477; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_479 = i == 10'h223 ? _GEN_478 : _GEN_477; // @[lut_mem_online.scala 247:34]
  wire  _GEN_480 = io_inputBit ? 1'h0 : _GEN_479; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_481 = i == 10'h223 ? _GEN_480 : _GEN_479; // @[lut_mem_online.scala 247:34]
  wire  _GEN_482 = ~io_inputBit ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_483 = i == 10'h224 ? _GEN_482 : _GEN_481; // @[lut_mem_online.scala 247:34]
  wire  _GEN_484 = io_inputBit | _GEN_483; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_485 = i == 10'h224 ? _GEN_484 : _GEN_483; // @[lut_mem_online.scala 247:34]
  wire  _GEN_486 = ~io_inputBit | _GEN_485; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_487 = i == 10'h225 ? _GEN_486 : _GEN_485; // @[lut_mem_online.scala 247:34]
  wire  _GEN_488 = io_inputBit ? 1'h0 : _GEN_487; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_489 = i == 10'h225 ? _GEN_488 : _GEN_487; // @[lut_mem_online.scala 247:34]
  wire  _GEN_490 = ~io_inputBit ? 1'h0 : _GEN_489; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_491 = i == 10'h226 ? _GEN_490 : _GEN_489; // @[lut_mem_online.scala 247:34]
  wire  _GEN_492 = io_inputBit | _GEN_491; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_493 = i == 10'h226 ? _GEN_492 : _GEN_491; // @[lut_mem_online.scala 247:34]
  wire  _GEN_494 = ~io_inputBit | _GEN_493; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_495 = i == 10'h227 ? _GEN_494 : _GEN_493; // @[lut_mem_online.scala 247:34]
  wire  _GEN_496 = io_inputBit ? 1'h0 : _GEN_495; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_497 = i == 10'h227 ? _GEN_496 : _GEN_495; // @[lut_mem_online.scala 247:34]
  wire  _GEN_498 = ~io_inputBit ? 1'h0 : _GEN_497; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_499 = i == 10'h228 ? _GEN_498 : _GEN_497; // @[lut_mem_online.scala 247:34]
  wire  _GEN_500 = io_inputBit | _GEN_499; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_501 = i == 10'h228 ? _GEN_500 : _GEN_499; // @[lut_mem_online.scala 247:34]
  wire  _GEN_502 = ~io_inputBit | _GEN_501; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_503 = i == 10'h229 ? _GEN_502 : _GEN_501; // @[lut_mem_online.scala 247:34]
  wire  _GEN_504 = io_inputBit ? 1'h0 : _GEN_503; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_505 = i == 10'h229 ? _GEN_504 : _GEN_503; // @[lut_mem_online.scala 247:34]
  wire  _GEN_506 = ~io_inputBit ? 1'h0 : _GEN_505; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_507 = i == 10'h22a ? _GEN_506 : _GEN_505; // @[lut_mem_online.scala 247:34]
  wire  _GEN_508 = io_inputBit | _GEN_507; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_509 = i == 10'h22a ? _GEN_508 : _GEN_507; // @[lut_mem_online.scala 247:34]
  wire  _GEN_510 = ~io_inputBit | _GEN_509; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_511 = i == 10'h22b ? _GEN_510 : _GEN_509; // @[lut_mem_online.scala 247:34]
  wire  _GEN_512 = io_inputBit ? 1'h0 : _GEN_511; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_513 = i == 10'h22b ? _GEN_512 : _GEN_511; // @[lut_mem_online.scala 247:34]
  wire  _GEN_514 = ~io_inputBit ? 1'h0 : _GEN_513; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_515 = i == 10'h22c ? _GEN_514 : _GEN_513; // @[lut_mem_online.scala 247:34]
  wire  _GEN_516 = io_inputBit | _GEN_515; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_517 = i == 10'h22c ? _GEN_516 : _GEN_515; // @[lut_mem_online.scala 247:34]
  wire  _GEN_518 = ~io_inputBit | _GEN_517; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_519 = i == 10'h22d ? _GEN_518 : _GEN_517; // @[lut_mem_online.scala 247:34]
  wire  _GEN_520 = io_inputBit ? 1'h0 : _GEN_519; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_521 = i == 10'h22d ? _GEN_520 : _GEN_519; // @[lut_mem_online.scala 247:34]
  wire  _GEN_522 = ~io_inputBit ? 1'h0 : _GEN_521; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_523 = i == 10'h22e ? _GEN_522 : _GEN_521; // @[lut_mem_online.scala 247:34]
  wire  _GEN_524 = io_inputBit | _GEN_523; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_525 = i == 10'h22e ? _GEN_524 : _GEN_523; // @[lut_mem_online.scala 247:34]
  wire  _GEN_526 = ~io_inputBit | _GEN_525; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_527 = i == 10'h22f ? _GEN_526 : _GEN_525; // @[lut_mem_online.scala 247:34]
  wire  _GEN_528 = io_inputBit ? 1'h0 : _GEN_527; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_529 = i == 10'h22f ? _GEN_528 : _GEN_527; // @[lut_mem_online.scala 247:34]
  wire  _GEN_530 = ~io_inputBit ? 1'h0 : _GEN_529; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_531 = i == 10'h230 ? _GEN_530 : _GEN_529; // @[lut_mem_online.scala 247:34]
  wire  _GEN_532 = io_inputBit | _GEN_531; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_533 = i == 10'h230 ? _GEN_532 : _GEN_531; // @[lut_mem_online.scala 247:34]
  wire  _GEN_534 = ~io_inputBit | _GEN_533; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_535 = i == 10'h231 ? _GEN_534 : _GEN_533; // @[lut_mem_online.scala 247:34]
  wire  _GEN_536 = io_inputBit ? 1'h0 : _GEN_535; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_537 = i == 10'h231 ? _GEN_536 : _GEN_535; // @[lut_mem_online.scala 247:34]
  wire  _GEN_538 = ~io_inputBit ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_539 = i == 10'h232 ? _GEN_538 : _GEN_537; // @[lut_mem_online.scala 247:34]
  wire  _GEN_540 = io_inputBit | _GEN_539; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_541 = i == 10'h232 ? _GEN_540 : _GEN_539; // @[lut_mem_online.scala 247:34]
  wire  _GEN_542 = ~io_inputBit | _GEN_541; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_543 = i == 10'h233 ? _GEN_542 : _GEN_541; // @[lut_mem_online.scala 247:34]
  wire  _GEN_544 = io_inputBit ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_545 = i == 10'h233 ? _GEN_544 : _GEN_543; // @[lut_mem_online.scala 247:34]
  wire  _GEN_546 = ~io_inputBit ? 1'h0 : _GEN_545; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_547 = i == 10'h234 ? _GEN_546 : _GEN_545; // @[lut_mem_online.scala 247:34]
  wire  _GEN_548 = io_inputBit | _GEN_547; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_549 = i == 10'h234 ? _GEN_548 : _GEN_547; // @[lut_mem_online.scala 247:34]
  wire  _GEN_550 = ~io_inputBit | _GEN_549; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_551 = i == 10'h235 ? _GEN_550 : _GEN_549; // @[lut_mem_online.scala 247:34]
  wire  _GEN_552 = io_inputBit ? 1'h0 : _GEN_551; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_553 = i == 10'h235 ? _GEN_552 : _GEN_551; // @[lut_mem_online.scala 247:34]
  wire  _GEN_554 = ~io_inputBit ? 1'h0 : _GEN_553; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_555 = i == 10'h236 ? _GEN_554 : _GEN_553; // @[lut_mem_online.scala 247:34]
  wire  _GEN_556 = io_inputBit | _GEN_555; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_557 = i == 10'h236 ? _GEN_556 : _GEN_555; // @[lut_mem_online.scala 247:34]
  wire  _GEN_558 = ~io_inputBit | _GEN_557; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_559 = i == 10'h237 ? _GEN_558 : _GEN_557; // @[lut_mem_online.scala 247:34]
  wire  _GEN_560 = io_inputBit ? 1'h0 : _GEN_559; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_561 = i == 10'h237 ? _GEN_560 : _GEN_559; // @[lut_mem_online.scala 247:34]
  wire  _GEN_562 = ~io_inputBit ? 1'h0 : _GEN_561; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_563 = i == 10'h238 ? _GEN_562 : _GEN_561; // @[lut_mem_online.scala 247:34]
  wire  _GEN_564 = io_inputBit | _GEN_563; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_565 = i == 10'h238 ? _GEN_564 : _GEN_563; // @[lut_mem_online.scala 247:34]
  wire  _GEN_566 = ~io_inputBit | _GEN_565; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_567 = i == 10'h239 ? _GEN_566 : _GEN_565; // @[lut_mem_online.scala 247:34]
  wire  _GEN_568 = io_inputBit ? 1'h0 : _GEN_567; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_569 = i == 10'h239 ? _GEN_568 : _GEN_567; // @[lut_mem_online.scala 247:34]
  wire  _GEN_570 = ~io_inputBit ? 1'h0 : _GEN_569; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_571 = i == 10'h23a ? _GEN_570 : _GEN_569; // @[lut_mem_online.scala 247:34]
  wire  _GEN_572 = io_inputBit | _GEN_571; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_573 = i == 10'h23a ? _GEN_572 : _GEN_571; // @[lut_mem_online.scala 247:34]
  wire  _GEN_574 = ~io_inputBit | _GEN_573; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_575 = i == 10'h23b ? _GEN_574 : _GEN_573; // @[lut_mem_online.scala 247:34]
  wire  _GEN_576 = io_inputBit ? 1'h0 : _GEN_575; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_577 = i == 10'h23b ? _GEN_576 : _GEN_575; // @[lut_mem_online.scala 247:34]
  wire  _GEN_578 = ~io_inputBit ? 1'h0 : _GEN_577; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_579 = i == 10'h23c ? _GEN_578 : _GEN_577; // @[lut_mem_online.scala 247:34]
  wire  _GEN_580 = io_inputBit | _GEN_579; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_581 = i == 10'h23c ? _GEN_580 : _GEN_579; // @[lut_mem_online.scala 247:34]
  wire  _GEN_582 = ~io_inputBit | _GEN_581; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_583 = i == 10'h23d ? _GEN_582 : _GEN_581; // @[lut_mem_online.scala 247:34]
  wire  _GEN_584 = io_inputBit ? 1'h0 : _GEN_583; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_585 = i == 10'h23d ? _GEN_584 : _GEN_583; // @[lut_mem_online.scala 247:34]
  wire  _GEN_586 = ~io_inputBit ? 1'h0 : _GEN_585; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_587 = i == 10'h23e ? _GEN_586 : _GEN_585; // @[lut_mem_online.scala 247:34]
  wire  _GEN_588 = io_inputBit | _GEN_587; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_589 = i == 10'h23e ? _GEN_588 : _GEN_587; // @[lut_mem_online.scala 247:34]
  wire  _GEN_590 = ~io_inputBit | _GEN_589; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_591 = i == 10'h23f ? _GEN_590 : _GEN_589; // @[lut_mem_online.scala 247:34]
  wire  _GEN_592 = io_inputBit ? 1'h0 : _GEN_591; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_593 = i == 10'h23f ? _GEN_592 : _GEN_591; // @[lut_mem_online.scala 247:34]
  wire  _GEN_594 = ~io_inputBit ? 1'h0 : _GEN_593; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_595 = i == 10'h240 ? _GEN_594 : _GEN_593; // @[lut_mem_online.scala 247:34]
  wire  _GEN_596 = io_inputBit | _GEN_595; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_597 = i == 10'h240 ? _GEN_596 : _GEN_595; // @[lut_mem_online.scala 247:34]
  wire  _GEN_598 = ~io_inputBit | _GEN_597; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_599 = i == 10'h241 ? _GEN_598 : _GEN_597; // @[lut_mem_online.scala 247:34]
  wire  _GEN_600 = io_inputBit ? 1'h0 : _GEN_599; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_601 = i == 10'h241 ? _GEN_600 : _GEN_599; // @[lut_mem_online.scala 247:34]
  wire  _GEN_602 = ~io_inputBit ? 1'h0 : _GEN_601; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_603 = i == 10'h242 ? _GEN_602 : _GEN_601; // @[lut_mem_online.scala 247:34]
  wire  _GEN_604 = io_inputBit | _GEN_603; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_605 = i == 10'h242 ? _GEN_604 : _GEN_603; // @[lut_mem_online.scala 247:34]
  wire  _GEN_606 = ~io_inputBit | _GEN_605; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_607 = i == 10'h243 ? _GEN_606 : _GEN_605; // @[lut_mem_online.scala 247:34]
  wire  _GEN_608 = io_inputBit ? 1'h0 : _GEN_607; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_609 = i == 10'h243 ? _GEN_608 : _GEN_607; // @[lut_mem_online.scala 247:34]
  wire  _GEN_610 = ~io_inputBit ? 1'h0 : _GEN_609; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_611 = i == 10'h244 ? _GEN_610 : _GEN_609; // @[lut_mem_online.scala 247:34]
  wire  _GEN_612 = io_inputBit | _GEN_611; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_613 = i == 10'h244 ? _GEN_612 : _GEN_611; // @[lut_mem_online.scala 247:34]
  wire  _GEN_614 = ~io_inputBit | _GEN_613; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_615 = i == 10'h245 ? _GEN_614 : _GEN_613; // @[lut_mem_online.scala 247:34]
  wire  _GEN_616 = io_inputBit ? 1'h0 : _GEN_615; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_617 = i == 10'h245 ? _GEN_616 : _GEN_615; // @[lut_mem_online.scala 247:34]
  wire  _GEN_618 = ~io_inputBit ? 1'h0 : _GEN_617; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_619 = i == 10'h246 ? _GEN_618 : _GEN_617; // @[lut_mem_online.scala 247:34]
  wire  _GEN_620 = io_inputBit | _GEN_619; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_621 = i == 10'h246 ? _GEN_620 : _GEN_619; // @[lut_mem_online.scala 247:34]
  wire  _GEN_622 = ~io_inputBit | _GEN_621; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_623 = i == 10'h247 ? _GEN_622 : _GEN_621; // @[lut_mem_online.scala 247:34]
  wire  _GEN_624 = io_inputBit ? 1'h0 : _GEN_623; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_625 = i == 10'h247 ? _GEN_624 : _GEN_623; // @[lut_mem_online.scala 247:34]
  wire  _GEN_626 = ~io_inputBit ? 1'h0 : _GEN_625; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_627 = i == 10'h248 ? _GEN_626 : _GEN_625; // @[lut_mem_online.scala 247:34]
  wire  _GEN_628 = io_inputBit | _GEN_627; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_629 = i == 10'h248 ? _GEN_628 : _GEN_627; // @[lut_mem_online.scala 247:34]
  wire  _GEN_630 = ~io_inputBit | _GEN_629; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_631 = i == 10'h249 ? _GEN_630 : _GEN_629; // @[lut_mem_online.scala 247:34]
  wire  _GEN_634 = io_inputBit ? 1'h0 : buffer_6; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_635 = i == 10'h0 ? _GEN_634 : buffer_6; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_636 = io_inputBit ? 1'h0 : _GEN_635; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_637 = i == 10'h1 ? _GEN_636 : _GEN_635; // @[lut_mem_online.scala 247:34]
  wire  _GEN_638 = io_inputBit ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_639 = i == 10'h8 ? _GEN_638 : _GEN_637; // @[lut_mem_online.scala 247:34]
  wire  _GEN_640 = ~io_inputBit ? 1'h0 : _GEN_639; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_641 = i == 10'hf ? _GEN_640 : _GEN_639; // @[lut_mem_online.scala 247:34]
  wire  _GEN_642 = io_inputBit ? 1'h0 : _GEN_641; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_643 = i == 10'h11 ? _GEN_642 : _GEN_641; // @[lut_mem_online.scala 247:34]
  wire  _GEN_644 = ~io_inputBit ? 1'h0 : _GEN_643; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_645 = i == 10'h20 ? _GEN_644 : _GEN_643; // @[lut_mem_online.scala 247:34]
  wire  _GEN_646 = io_inputBit ? 1'h0 : _GEN_645; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_647 = i == 10'h48 ? _GEN_646 : _GEN_645; // @[lut_mem_online.scala 247:34]
  wire  _GEN_648 = ~io_inputBit ? 1'h0 : _GEN_647; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_649 = i == 10'h10b ? _GEN_648 : _GEN_647; // @[lut_mem_online.scala 247:34]
  wire  _GEN_650 = io_inputBit ? 1'h0 : _GEN_649; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_651 = i == 10'h124 ? _GEN_650 : _GEN_649; // @[lut_mem_online.scala 247:34]
  wire  _GEN_652 = ~io_inputBit ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_653 = i == 10'h218 ? _GEN_652 : _GEN_651; // @[lut_mem_online.scala 247:34]
  wire  _GEN_654 = io_inputBit | _GEN_653; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_655 = i == 10'h218 ? _GEN_654 : _GEN_653; // @[lut_mem_online.scala 247:34]
  wire  _GEN_656 = ~io_inputBit ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_657 = i == 10'h219 ? _GEN_656 : _GEN_655; // @[lut_mem_online.scala 247:34]
  wire  _GEN_658 = io_inputBit | _GEN_657; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_659 = i == 10'h219 ? _GEN_658 : _GEN_657; // @[lut_mem_online.scala 247:34]
  wire  _GEN_660 = ~io_inputBit ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_661 = i == 10'h21a ? _GEN_660 : _GEN_659; // @[lut_mem_online.scala 247:34]
  wire  _GEN_662 = io_inputBit | _GEN_661; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_663 = i == 10'h21a ? _GEN_662 : _GEN_661; // @[lut_mem_online.scala 247:34]
  wire  _GEN_664 = ~io_inputBit ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_665 = i == 10'h21b ? _GEN_664 : _GEN_663; // @[lut_mem_online.scala 247:34]
  wire  _GEN_666 = io_inputBit | _GEN_665; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_667 = i == 10'h21b ? _GEN_666 : _GEN_665; // @[lut_mem_online.scala 247:34]
  wire  _GEN_668 = ~io_inputBit ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_669 = i == 10'h21c ? _GEN_668 : _GEN_667; // @[lut_mem_online.scala 247:34]
  wire  _GEN_670 = io_inputBit | _GEN_669; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_671 = i == 10'h21c ? _GEN_670 : _GEN_669; // @[lut_mem_online.scala 247:34]
  wire  _GEN_672 = ~io_inputBit ? 1'h0 : _GEN_671; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_673 = i == 10'h21d ? _GEN_672 : _GEN_671; // @[lut_mem_online.scala 247:34]
  wire  _GEN_674 = io_inputBit | _GEN_673; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_675 = i == 10'h21d ? _GEN_674 : _GEN_673; // @[lut_mem_online.scala 247:34]
  wire  _GEN_676 = ~io_inputBit ? 1'h0 : _GEN_675; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_677 = i == 10'h21e ? _GEN_676 : _GEN_675; // @[lut_mem_online.scala 247:34]
  wire  _GEN_678 = io_inputBit | _GEN_677; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_679 = i == 10'h21e ? _GEN_678 : _GEN_677; // @[lut_mem_online.scala 247:34]
  wire  _GEN_680 = ~io_inputBit ? 1'h0 : _GEN_679; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_681 = i == 10'h21f ? _GEN_680 : _GEN_679; // @[lut_mem_online.scala 247:34]
  wire  _GEN_682 = io_inputBit | _GEN_681; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_683 = i == 10'h21f ? _GEN_682 : _GEN_681; // @[lut_mem_online.scala 247:34]
  wire  _GEN_684 = ~io_inputBit ? 1'h0 : _GEN_683; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_685 = i == 10'h220 ? _GEN_684 : _GEN_683; // @[lut_mem_online.scala 247:34]
  wire  _GEN_686 = io_inputBit | _GEN_685; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_687 = i == 10'h220 ? _GEN_686 : _GEN_685; // @[lut_mem_online.scala 247:34]
  wire  _GEN_688 = ~io_inputBit ? 1'h0 : _GEN_687; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_689 = i == 10'h221 ? _GEN_688 : _GEN_687; // @[lut_mem_online.scala 247:34]
  wire  _GEN_690 = io_inputBit | _GEN_689; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_691 = i == 10'h221 ? _GEN_690 : _GEN_689; // @[lut_mem_online.scala 247:34]
  wire  _GEN_692 = ~io_inputBit ? 1'h0 : _GEN_691; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_693 = i == 10'h222 ? _GEN_692 : _GEN_691; // @[lut_mem_online.scala 247:34]
  wire  _GEN_694 = io_inputBit | _GEN_693; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_695 = i == 10'h222 ? _GEN_694 : _GEN_693; // @[lut_mem_online.scala 247:34]
  wire  _GEN_696 = ~io_inputBit ? 1'h0 : _GEN_695; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_697 = i == 10'h223 ? _GEN_696 : _GEN_695; // @[lut_mem_online.scala 247:34]
  wire  _GEN_698 = io_inputBit | _GEN_697; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_699 = i == 10'h223 ? _GEN_698 : _GEN_697; // @[lut_mem_online.scala 247:34]
  wire  _GEN_700 = ~io_inputBit ? 1'h0 : _GEN_699; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_701 = i == 10'h224 ? _GEN_700 : _GEN_699; // @[lut_mem_online.scala 247:34]
  wire  _GEN_702 = io_inputBit | _GEN_701; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_703 = i == 10'h224 ? _GEN_702 : _GEN_701; // @[lut_mem_online.scala 247:34]
  wire  _GEN_704 = ~io_inputBit ? 1'h0 : _GEN_703; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_705 = i == 10'h225 ? _GEN_704 : _GEN_703; // @[lut_mem_online.scala 247:34]
  wire  _GEN_706 = io_inputBit | _GEN_705; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_707 = i == 10'h225 ? _GEN_706 : _GEN_705; // @[lut_mem_online.scala 247:34]
  wire  _GEN_708 = ~io_inputBit ? 1'h0 : _GEN_707; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_709 = i == 10'h226 ? _GEN_708 : _GEN_707; // @[lut_mem_online.scala 247:34]
  wire  _GEN_710 = io_inputBit | _GEN_709; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_711 = i == 10'h226 ? _GEN_710 : _GEN_709; // @[lut_mem_online.scala 247:34]
  wire  _GEN_712 = ~io_inputBit ? 1'h0 : _GEN_711; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_713 = i == 10'h227 ? _GEN_712 : _GEN_711; // @[lut_mem_online.scala 247:34]
  wire  _GEN_714 = io_inputBit | _GEN_713; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_715 = i == 10'h227 ? _GEN_714 : _GEN_713; // @[lut_mem_online.scala 247:34]
  wire  _GEN_716 = ~io_inputBit ? 1'h0 : _GEN_715; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_717 = i == 10'h228 ? _GEN_716 : _GEN_715; // @[lut_mem_online.scala 247:34]
  wire  _GEN_718 = io_inputBit | _GEN_717; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_719 = i == 10'h228 ? _GEN_718 : _GEN_717; // @[lut_mem_online.scala 247:34]
  wire  _GEN_720 = ~io_inputBit ? 1'h0 : _GEN_719; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_721 = i == 10'h229 ? _GEN_720 : _GEN_719; // @[lut_mem_online.scala 247:34]
  wire  _GEN_722 = io_inputBit | _GEN_721; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_723 = i == 10'h229 ? _GEN_722 : _GEN_721; // @[lut_mem_online.scala 247:34]
  wire  _GEN_724 = ~io_inputBit ? 1'h0 : _GEN_723; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_725 = i == 10'h22a ? _GEN_724 : _GEN_723; // @[lut_mem_online.scala 247:34]
  wire  _GEN_726 = io_inputBit | _GEN_725; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_727 = i == 10'h22a ? _GEN_726 : _GEN_725; // @[lut_mem_online.scala 247:34]
  wire  _GEN_728 = ~io_inputBit ? 1'h0 : _GEN_727; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_729 = i == 10'h22b ? _GEN_728 : _GEN_727; // @[lut_mem_online.scala 247:34]
  wire  _GEN_730 = io_inputBit | _GEN_729; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_731 = i == 10'h22b ? _GEN_730 : _GEN_729; // @[lut_mem_online.scala 247:34]
  wire  _GEN_732 = ~io_inputBit ? 1'h0 : _GEN_731; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_733 = i == 10'h22c ? _GEN_732 : _GEN_731; // @[lut_mem_online.scala 247:34]
  wire  _GEN_734 = io_inputBit | _GEN_733; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_735 = i == 10'h22c ? _GEN_734 : _GEN_733; // @[lut_mem_online.scala 247:34]
  wire  _GEN_736 = ~io_inputBit ? 1'h0 : _GEN_735; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_737 = i == 10'h22d ? _GEN_736 : _GEN_735; // @[lut_mem_online.scala 247:34]
  wire  _GEN_738 = io_inputBit | _GEN_737; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_739 = i == 10'h22d ? _GEN_738 : _GEN_737; // @[lut_mem_online.scala 247:34]
  wire  _GEN_740 = ~io_inputBit ? 1'h0 : _GEN_739; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_741 = i == 10'h22e ? _GEN_740 : _GEN_739; // @[lut_mem_online.scala 247:34]
  wire  _GEN_742 = io_inputBit | _GEN_741; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_743 = i == 10'h22e ? _GEN_742 : _GEN_741; // @[lut_mem_online.scala 247:34]
  wire  _GEN_744 = ~io_inputBit ? 1'h0 : _GEN_743; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_745 = i == 10'h22f ? _GEN_744 : _GEN_743; // @[lut_mem_online.scala 247:34]
  wire  _GEN_746 = io_inputBit | _GEN_745; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_747 = i == 10'h22f ? _GEN_746 : _GEN_745; // @[lut_mem_online.scala 247:34]
  wire  _GEN_748 = ~io_inputBit ? 1'h0 : _GEN_747; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_749 = i == 10'h230 ? _GEN_748 : _GEN_747; // @[lut_mem_online.scala 247:34]
  wire  _GEN_750 = io_inputBit | _GEN_749; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_751 = i == 10'h230 ? _GEN_750 : _GEN_749; // @[lut_mem_online.scala 247:34]
  wire  _GEN_752 = ~io_inputBit ? 1'h0 : _GEN_751; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_753 = i == 10'h231 ? _GEN_752 : _GEN_751; // @[lut_mem_online.scala 247:34]
  wire  _GEN_754 = io_inputBit | _GEN_753; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_755 = i == 10'h231 ? _GEN_754 : _GEN_753; // @[lut_mem_online.scala 247:34]
  wire  _GEN_756 = ~io_inputBit ? 1'h0 : _GEN_755; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_757 = i == 10'h232 ? _GEN_756 : _GEN_755; // @[lut_mem_online.scala 247:34]
  wire  _GEN_758 = io_inputBit | _GEN_757; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_759 = i == 10'h232 ? _GEN_758 : _GEN_757; // @[lut_mem_online.scala 247:34]
  wire  _GEN_760 = ~io_inputBit ? 1'h0 : _GEN_759; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_761 = i == 10'h233 ? _GEN_760 : _GEN_759; // @[lut_mem_online.scala 247:34]
  wire  _GEN_762 = io_inputBit | _GEN_761; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_763 = i == 10'h233 ? _GEN_762 : _GEN_761; // @[lut_mem_online.scala 247:34]
  wire  _GEN_764 = ~io_inputBit ? 1'h0 : _GEN_763; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_765 = i == 10'h234 ? _GEN_764 : _GEN_763; // @[lut_mem_online.scala 247:34]
  wire  _GEN_766 = io_inputBit | _GEN_765; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_767 = i == 10'h234 ? _GEN_766 : _GEN_765; // @[lut_mem_online.scala 247:34]
  wire  _GEN_768 = ~io_inputBit ? 1'h0 : _GEN_767; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_769 = i == 10'h235 ? _GEN_768 : _GEN_767; // @[lut_mem_online.scala 247:34]
  wire  _GEN_770 = io_inputBit | _GEN_769; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_771 = i == 10'h235 ? _GEN_770 : _GEN_769; // @[lut_mem_online.scala 247:34]
  wire  _GEN_772 = ~io_inputBit ? 1'h0 : _GEN_771; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_773 = i == 10'h236 ? _GEN_772 : _GEN_771; // @[lut_mem_online.scala 247:34]
  wire  _GEN_774 = io_inputBit | _GEN_773; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_775 = i == 10'h236 ? _GEN_774 : _GEN_773; // @[lut_mem_online.scala 247:34]
  wire  _GEN_776 = ~io_inputBit ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_777 = i == 10'h237 ? _GEN_776 : _GEN_775; // @[lut_mem_online.scala 247:34]
  wire  _GEN_778 = io_inputBit | _GEN_777; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_779 = i == 10'h237 ? _GEN_778 : _GEN_777; // @[lut_mem_online.scala 247:34]
  wire  _GEN_780 = ~io_inputBit ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_781 = i == 10'h238 ? _GEN_780 : _GEN_779; // @[lut_mem_online.scala 247:34]
  wire  _GEN_782 = io_inputBit | _GEN_781; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_783 = i == 10'h238 ? _GEN_782 : _GEN_781; // @[lut_mem_online.scala 247:34]
  wire  _GEN_784 = ~io_inputBit ? 1'h0 : _GEN_783; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_785 = i == 10'h239 ? _GEN_784 : _GEN_783; // @[lut_mem_online.scala 247:34]
  wire  _GEN_786 = io_inputBit | _GEN_785; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_787 = i == 10'h239 ? _GEN_786 : _GEN_785; // @[lut_mem_online.scala 247:34]
  wire  _GEN_788 = ~io_inputBit ? 1'h0 : _GEN_787; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_789 = i == 10'h23a ? _GEN_788 : _GEN_787; // @[lut_mem_online.scala 247:34]
  wire  _GEN_790 = io_inputBit | _GEN_789; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_791 = i == 10'h23a ? _GEN_790 : _GEN_789; // @[lut_mem_online.scala 247:34]
  wire  _GEN_792 = ~io_inputBit ? 1'h0 : _GEN_791; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_793 = i == 10'h23b ? _GEN_792 : _GEN_791; // @[lut_mem_online.scala 247:34]
  wire  _GEN_794 = io_inputBit | _GEN_793; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_795 = i == 10'h23b ? _GEN_794 : _GEN_793; // @[lut_mem_online.scala 247:34]
  wire  _GEN_796 = ~io_inputBit ? 1'h0 : _GEN_795; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_797 = i == 10'h23c ? _GEN_796 : _GEN_795; // @[lut_mem_online.scala 247:34]
  wire  _GEN_798 = io_inputBit | _GEN_797; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_799 = i == 10'h23c ? _GEN_798 : _GEN_797; // @[lut_mem_online.scala 247:34]
  wire  _GEN_800 = ~io_inputBit ? 1'h0 : _GEN_799; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_801 = i == 10'h23d ? _GEN_800 : _GEN_799; // @[lut_mem_online.scala 247:34]
  wire  _GEN_802 = io_inputBit | _GEN_801; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_803 = i == 10'h23d ? _GEN_802 : _GEN_801; // @[lut_mem_online.scala 247:34]
  wire  _GEN_804 = ~io_inputBit ? 1'h0 : _GEN_803; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_805 = i == 10'h23e ? _GEN_804 : _GEN_803; // @[lut_mem_online.scala 247:34]
  wire  _GEN_806 = io_inputBit | _GEN_805; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_807 = i == 10'h23e ? _GEN_806 : _GEN_805; // @[lut_mem_online.scala 247:34]
  wire  _GEN_808 = ~io_inputBit ? 1'h0 : _GEN_807; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_809 = i == 10'h23f ? _GEN_808 : _GEN_807; // @[lut_mem_online.scala 247:34]
  wire  _GEN_810 = io_inputBit | _GEN_809; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_811 = i == 10'h23f ? _GEN_810 : _GEN_809; // @[lut_mem_online.scala 247:34]
  wire  _GEN_812 = ~io_inputBit ? 1'h0 : _GEN_811; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_813 = i == 10'h240 ? _GEN_812 : _GEN_811; // @[lut_mem_online.scala 247:34]
  wire  _GEN_814 = io_inputBit | _GEN_813; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_815 = i == 10'h240 ? _GEN_814 : _GEN_813; // @[lut_mem_online.scala 247:34]
  wire  _GEN_816 = ~io_inputBit ? 1'h0 : _GEN_815; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_817 = i == 10'h241 ? _GEN_816 : _GEN_815; // @[lut_mem_online.scala 247:34]
  wire  _GEN_818 = io_inputBit | _GEN_817; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_819 = i == 10'h241 ? _GEN_818 : _GEN_817; // @[lut_mem_online.scala 247:34]
  wire  _GEN_820 = ~io_inputBit ? 1'h0 : _GEN_819; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_821 = i == 10'h242 ? _GEN_820 : _GEN_819; // @[lut_mem_online.scala 247:34]
  wire  _GEN_822 = io_inputBit | _GEN_821; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_823 = i == 10'h242 ? _GEN_822 : _GEN_821; // @[lut_mem_online.scala 247:34]
  wire  _GEN_824 = ~io_inputBit ? 1'h0 : _GEN_823; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_825 = i == 10'h243 ? _GEN_824 : _GEN_823; // @[lut_mem_online.scala 247:34]
  wire  _GEN_826 = io_inputBit | _GEN_825; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_827 = i == 10'h243 ? _GEN_826 : _GEN_825; // @[lut_mem_online.scala 247:34]
  wire  _GEN_828 = ~io_inputBit ? 1'h0 : _GEN_827; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_829 = i == 10'h244 ? _GEN_828 : _GEN_827; // @[lut_mem_online.scala 247:34]
  wire  _GEN_830 = io_inputBit | _GEN_829; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_831 = i == 10'h244 ? _GEN_830 : _GEN_829; // @[lut_mem_online.scala 247:34]
  wire  _GEN_832 = ~io_inputBit ? 1'h0 : _GEN_831; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_833 = i == 10'h245 ? _GEN_832 : _GEN_831; // @[lut_mem_online.scala 247:34]
  wire  _GEN_834 = io_inputBit | _GEN_833; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_835 = i == 10'h245 ? _GEN_834 : _GEN_833; // @[lut_mem_online.scala 247:34]
  wire  _GEN_836 = ~io_inputBit ? 1'h0 : _GEN_835; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_837 = i == 10'h246 ? _GEN_836 : _GEN_835; // @[lut_mem_online.scala 247:34]
  wire  _GEN_838 = io_inputBit | _GEN_837; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_839 = i == 10'h246 ? _GEN_838 : _GEN_837; // @[lut_mem_online.scala 247:34]
  wire  _GEN_840 = ~io_inputBit ? 1'h0 : _GEN_839; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_841 = i == 10'h247 ? _GEN_840 : _GEN_839; // @[lut_mem_online.scala 247:34]
  wire  _GEN_842 = io_inputBit | _GEN_841; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_843 = i == 10'h247 ? _GEN_842 : _GEN_841; // @[lut_mem_online.scala 247:34]
  wire  _GEN_844 = ~io_inputBit ? 1'h0 : _GEN_843; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_845 = i == 10'h248 ? _GEN_844 : _GEN_843; // @[lut_mem_online.scala 247:34]
  wire  _GEN_846 = io_inputBit | _GEN_845; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_847 = i == 10'h248 ? _GEN_846 : _GEN_845; // @[lut_mem_online.scala 247:34]
  wire  _GEN_848 = ~io_inputBit ? 1'h0 : _GEN_847; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_849 = i == 10'h249 ? _GEN_848 : _GEN_847; // @[lut_mem_online.scala 247:34]
  wire  _GEN_850 = io_inputBit | _GEN_849; // @[lut_mem_online.scala 249:46 251:32]
  wire  _T_855 = counter < 5'h11; // @[lut_mem_online.scala 262:22]
  wire  _T_857 = counter >= 5'ha; // @[lut_mem_online.scala 270:30]
  wire [4:0] _outResult_T_1 = counter - 5'ha; // @[lut_mem_online.scala 272:41]
  wire  _GEN_860 = 4'h1 == _outResult_T_1[3:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_861 = 4'h2 == _outResult_T_1[3:0] ? buffer_2 : _GEN_860; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_862 = 4'h3 == _outResult_T_1[3:0] ? buffer_3 : _GEN_861; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_863 = 4'h4 == _outResult_T_1[3:0] ? buffer_4 : _GEN_862; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_864 = 4'h5 == _outResult_T_1[3:0] ? buffer_5 : _GEN_863; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_865 = 4'h6 == _outResult_T_1[3:0] ? buffer_6 : _GEN_864; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_866 = 4'h7 == _outResult_T_1[3:0] ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_867 = 4'h8 == _outResult_T_1[3:0] ? 1'h0 : _GEN_866; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_868 = 4'h9 == _outResult_T_1[3:0] ? 1'h0 : _GEN_867; // @[lut_mem_online.scala 272:{23,23}]
  wire  _T_861 = ~reset; // @[lut_mem_online.scala 278:21]
  wire  _GEN_870 = counter >= 5'ha ? _GEN_868 : outResult; // @[lut_mem_online.scala 270:42 272:23 224:26]
  wire  _GEN_872 = _T_2 ? 1'h0 : _GEN_870; // @[lut_mem_online.scala 267:35 269:23]
  wire  _T_862 = i < 10'h1ff; // @[lut_mem_online.scala 293:18]
  wire [11:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 307:24]
  wire [11:0] _i_T_2 = _i_T + 12'h1; // @[lut_mem_online.scala 307:28]
  wire [11:0] _i_T_5 = _i_T + 12'h2; // @[lut_mem_online.scala 309:28]
  wire [11:0] _GEN_873 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 308:45 309:17 215:18]
  wire [11:0] _GEN_874 = _T_10 ? _i_T_2 : _GEN_873; // @[lut_mem_online.scala 306:39 307:17]
  wire  _T_867 = i < 10'h3ff; // @[lut_mem_online.scala 316:24]
  wire [9:0] _GEN_875 = i < 10'h3ff ? 10'h3ff : i; // @[lut_mem_online.scala 316:63 324:15 215:18]
  wire [11:0] _GEN_876 = i < 10'h1ff ? _GEN_874 : {{2'd0}, _GEN_875}; // @[lut_mem_online.scala 293:61]
  wire [4:0] _counter_T_1 = counter + 5'h1; // @[lut_mem_online.scala 327:30]
  wire  _GEN_878 = counter < 5'h11 & _GEN_872; // @[lut_mem_online.scala 262:52 335:21]
  wire [11:0] _GEN_879 = counter < 5'h11 ? _GEN_876 : {{2'd0}, i}; // @[lut_mem_online.scala 215:18 262:52]
  wire  _GEN_902 = io_start & _GEN_878; // @[lut_mem_online.scala 229:29 362:15]
  wire [11:0] _GEN_903 = io_start ? _GEN_879 : 12'h0; // @[lut_mem_online.scala 229:29 360:7]
  wire [11:0] _GEN_906 = reset ? 12'h0 : _GEN_903; // @[lut_mem_online.scala 215:{18,18}]
  wire  _GEN_907 = io_start & _T_855; // @[lut_mem_online.scala 278:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 369:16]
  always @(posedge clock) begin
    i <= _GEN_906[9:0]; // @[lut_mem_online.scala 215:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h22a) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_0 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_0 <= _GEN_19;
          end
        end else begin
          buffer_0 <= _GEN_19;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h23a) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_1 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_1 <= _GEN_63;
          end
        end else begin
          buffer_1 <= _GEN_63;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h242) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_2 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_2 <= _GEN_137;
          end
        end else begin
          buffer_2 <= _GEN_137;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h246) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_3 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_3 <= _GEN_247;
          end
        end else begin
          buffer_3 <= _GEN_247;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h248) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_4 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_4 <= _GEN_413;
          end
        end else begin
          buffer_4 <= _GEN_413;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h249) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_5 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_5 <= _GEN_631;
          end
        end else begin
          buffer_5 <= _GEN_631;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h249) begin // @[lut_mem_online.scala 247:34]
          buffer_6 <= _GEN_850;
        end else if (i == 10'h249) begin // @[lut_mem_online.scala 247:34]
          buffer_6 <= _GEN_848;
        end else begin
          buffer_6 <= _GEN_847;
        end
      end
    end
    if (reset) begin // @[lut_mem_online.scala 221:24]
      counter <= 5'h0; // @[lut_mem_online.scala 221:24]
    end else if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'h11) begin // @[lut_mem_online.scala 262:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 327:19]
      end
    end else begin
      counter <= 5'h0; // @[lut_mem_online.scala 361:13]
    end
    if (reset) begin // @[lut_mem_online.scala 224:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 224:26]
    end else begin
      outResult <= _GEN_902;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_855 & ~_T_2 & _T_857 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 278:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_907 & _T_862 & _T_861) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 300:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_907 & ~_T_862 & _T_867 & _T_861) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 319:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
