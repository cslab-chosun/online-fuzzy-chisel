module LutMembershipFunctionOnline_7(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [7:0] i; // @[lut_mem_online.scala 206:18]
  reg  buffer_0; // @[lut_mem_online.scala 210:19]
  reg  buffer_1; // @[lut_mem_online.scala 210:19]
  reg  buffer_2; // @[lut_mem_online.scala 210:19]
  reg  buffer_3; // @[lut_mem_online.scala 210:19]
  reg  buffer_4; // @[lut_mem_online.scala 210:19]
  reg  buffer_5; // @[lut_mem_online.scala 210:19]
  reg  buffer_6; // @[lut_mem_online.scala 210:19]
  reg [4:0] counter; // @[lut_mem_online.scala 212:24]
  reg  outResult; // @[lut_mem_online.scala 215:26]
  wire  _GEN_0 = io_inputBit ? 1'h0 : buffer_0; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_1 = i == 8'h0 ? _GEN_0 : buffer_0; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_2 = io_inputBit ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3 = i == 8'h1 ? _GEN_2 : _GEN_1; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4 = io_inputBit ? 1'h0 : _GEN_3; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5 = i == 8'h3 ? _GEN_4 : _GEN_3; // @[lut_mem_online.scala 235:34]
  wire  _T_10 = ~io_inputBit; // @[lut_mem_online.scala 237:32]
  wire  _GEN_6 = ~io_inputBit | _GEN_5; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_7 = i == 8'h7 ? _GEN_6 : _GEN_5; // @[lut_mem_online.scala 235:34]
  wire  _GEN_8 = io_inputBit ? 1'h0 : _GEN_7; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_9 = i == 8'h10 ? _GEN_8 : _GEN_7; // @[lut_mem_online.scala 235:34]
  wire  _GEN_10 = ~io_inputBit | _GEN_9; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_11 = i == 8'h21 ? _GEN_10 : _GEN_9; // @[lut_mem_online.scala 235:34]
  wire  _GEN_12 = io_inputBit ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_13 = i == 8'h44 ? _GEN_12 : _GEN_11; // @[lut_mem_online.scala 235:34]
  wire  _GEN_14 = ~io_inputBit | _GEN_13; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_15 = i == 8'h89 ? _GEN_14 : _GEN_13; // @[lut_mem_online.scala 235:34]
  wire [8:0] _GEN_6084 = {{1'd0}, i}; // @[lut_mem_online.scala 235:20]
  wire  _GEN_16 = ~io_inputBit | _GEN_15; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_17 = _GEN_6084 == 9'h114 ? _GEN_16 : _GEN_15; // @[lut_mem_online.scala 235:34]
  wire [9:0] _GEN_6085 = {{2'd0}, i}; // @[lut_mem_online.scala 235:20]
  wire  _GEN_18 = ~io_inputBit | _GEN_17; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_19 = _GEN_6085 == 10'h22a ? _GEN_18 : _GEN_17; // @[lut_mem_online.scala 235:34]
  wire  _GEN_20 = io_inputBit ? 1'h0 : _GEN_19; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_21 = _GEN_6085 == 10'h22a ? _GEN_20 : _GEN_19; // @[lut_mem_online.scala 235:34]
  wire  _GEN_22 = io_inputBit ? 1'h0 : buffer_1; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_23 = i == 8'h0 ? _GEN_22 : buffer_1; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_24 = io_inputBit ? 1'h0 : _GEN_23; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_25 = i == 8'h1 ? _GEN_24 : _GEN_23; // @[lut_mem_online.scala 235:34]
  wire  _GEN_26 = io_inputBit ? 1'h0 : _GEN_25; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_27 = i == 8'h3 ? _GEN_26 : _GEN_25; // @[lut_mem_online.scala 235:34]
  wire  _GEN_28 = ~io_inputBit | _GEN_27; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_29 = i == 8'hf ? _GEN_28 : _GEN_27; // @[lut_mem_online.scala 235:34]
  wire  _GEN_30 = ~io_inputBit | _GEN_29; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_31 = i == 8'h20 ? _GEN_30 : _GEN_29; // @[lut_mem_online.scala 235:34]
  wire  _GEN_32 = ~io_inputBit ? 1'h0 : _GEN_31; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_33 = i == 8'h21 ? _GEN_32 : _GEN_31; // @[lut_mem_online.scala 235:34]
  wire  _GEN_34 = ~io_inputBit | _GEN_33; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_35 = i == 8'h22 ? _GEN_34 : _GEN_33; // @[lut_mem_online.scala 235:34]
  wire  _GEN_36 = io_inputBit ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_37 = i == 8'h42 ? _GEN_36 : _GEN_35; // @[lut_mem_online.scala 235:34]
  wire  _GEN_38 = io_inputBit | _GEN_37; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_39 = i == 8'h44 ? _GEN_38 : _GEN_37; // @[lut_mem_online.scala 235:34]
  wire  _GEN_40 = io_inputBit ? 1'h0 : _GEN_39; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_41 = i == 8'h46 ? _GEN_40 : _GEN_39; // @[lut_mem_online.scala 235:34]
  wire  _GEN_42 = ~io_inputBit | _GEN_41; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_43 = i == 8'h85 ? _GEN_42 : _GEN_41; // @[lut_mem_online.scala 235:34]
  wire  _GEN_44 = ~io_inputBit ? 1'h0 : _GEN_43; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_45 = i == 8'h89 ? _GEN_44 : _GEN_43; // @[lut_mem_online.scala 235:34]
  wire  _GEN_46 = ~io_inputBit | _GEN_45; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_47 = i == 8'h8d ? _GEN_46 : _GEN_45; // @[lut_mem_online.scala 235:34]
  wire  _GEN_48 = ~io_inputBit | _GEN_47; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_49 = _GEN_6084 == 9'h10c ? _GEN_48 : _GEN_47; // @[lut_mem_online.scala 235:34]
  wire  _GEN_50 = ~io_inputBit ? 1'h0 : _GEN_49; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_51 = _GEN_6084 == 9'h114 ? _GEN_50 : _GEN_49; // @[lut_mem_online.scala 235:34]
  wire  _GEN_52 = ~io_inputBit | _GEN_51; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_53 = _GEN_6084 == 9'h11c ? _GEN_52 : _GEN_51; // @[lut_mem_online.scala 235:34]
  wire  _GEN_54 = ~io_inputBit | _GEN_53; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_55 = _GEN_6085 == 10'h21a ? _GEN_54 : _GEN_53; // @[lut_mem_online.scala 235:34]
  wire  _GEN_56 = io_inputBit ? 1'h0 : _GEN_55; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_57 = _GEN_6085 == 10'h21a ? _GEN_56 : _GEN_55; // @[lut_mem_online.scala 235:34]
  wire  _GEN_58 = ~io_inputBit ? 1'h0 : _GEN_57; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_59 = _GEN_6085 == 10'h22a ? _GEN_58 : _GEN_57; // @[lut_mem_online.scala 235:34]
  wire  _GEN_60 = io_inputBit | _GEN_59; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_61 = _GEN_6085 == 10'h22a ? _GEN_60 : _GEN_59; // @[lut_mem_online.scala 235:34]
  wire  _GEN_62 = ~io_inputBit | _GEN_61; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_63 = _GEN_6085 == 10'h23a ? _GEN_62 : _GEN_61; // @[lut_mem_online.scala 235:34]
  wire  _GEN_64 = io_inputBit ? 1'h0 : _GEN_63; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_65 = _GEN_6085 == 10'h23a ? _GEN_64 : _GEN_63; // @[lut_mem_online.scala 235:34]
  wire  _GEN_66 = io_inputBit ? 1'h0 : buffer_2; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_67 = i == 8'h0 ? _GEN_66 : buffer_2; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_68 = io_inputBit ? 1'h0 : _GEN_67; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_69 = i == 8'h1 ? _GEN_68 : _GEN_67; // @[lut_mem_online.scala 235:34]
  wire  _GEN_70 = io_inputBit ? 1'h0 : _GEN_69; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_71 = i == 8'h8 ? _GEN_70 : _GEN_69; // @[lut_mem_online.scala 235:34]
  wire  _GEN_72 = ~io_inputBit ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_73 = i == 8'hf ? _GEN_72 : _GEN_71; // @[lut_mem_online.scala 235:34]
  wire  _GEN_74 = io_inputBit ? 1'h0 : _GEN_73; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_75 = i == 8'h11 ? _GEN_74 : _GEN_73; // @[lut_mem_online.scala 235:34]
  wire  _GEN_76 = ~io_inputBit ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_77 = i == 8'h20 ? _GEN_76 : _GEN_75; // @[lut_mem_online.scala 235:34]
  wire  _GEN_78 = io_inputBit ? 1'h0 : _GEN_77; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_79 = i == 8'h23 ? _GEN_78 : _GEN_77; // @[lut_mem_online.scala 235:34]
  wire  _GEN_80 = io_inputBit | _GEN_79; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_81 = i == 8'h42 ? _GEN_80 : _GEN_79; // @[lut_mem_online.scala 235:34]
  wire  _GEN_82 = io_inputBit ? 1'h0 : _GEN_81; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_83 = i == 8'h43 ? _GEN_82 : _GEN_81; // @[lut_mem_online.scala 235:34]
  wire  _GEN_84 = io_inputBit | _GEN_83; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_85 = i == 8'h44 ? _GEN_84 : _GEN_83; // @[lut_mem_online.scala 235:34]
  wire  _GEN_86 = io_inputBit ? 1'h0 : _GEN_85; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_87 = i == 8'h45 ? _GEN_86 : _GEN_85; // @[lut_mem_online.scala 235:34]
  wire  _GEN_88 = io_inputBit | _GEN_87; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_89 = i == 8'h46 ? _GEN_88 : _GEN_87; // @[lut_mem_online.scala 235:34]
  wire  _GEN_90 = io_inputBit ? 1'h0 : _GEN_89; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_91 = i == 8'h47 ? _GEN_90 : _GEN_89; // @[lut_mem_online.scala 235:34]
  wire  _GEN_92 = ~io_inputBit ? 1'h0 : _GEN_91; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_93 = i == 8'h85 ? _GEN_92 : _GEN_91; // @[lut_mem_online.scala 235:34]
  wire  _GEN_94 = ~io_inputBit | _GEN_93; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_95 = i == 8'h87 ? _GEN_94 : _GEN_93; // @[lut_mem_online.scala 235:34]
  wire  _GEN_96 = ~io_inputBit ? 1'h0 : _GEN_95; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_97 = i == 8'h89 ? _GEN_96 : _GEN_95; // @[lut_mem_online.scala 235:34]
  wire  _GEN_98 = ~io_inputBit | _GEN_97; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_99 = i == 8'h8b ? _GEN_98 : _GEN_97; // @[lut_mem_online.scala 235:34]
  wire  _GEN_100 = ~io_inputBit ? 1'h0 : _GEN_99; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_101 = i == 8'h8d ? _GEN_100 : _GEN_99; // @[lut_mem_online.scala 235:34]
  wire  _GEN_102 = ~io_inputBit | _GEN_101; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_103 = i == 8'h8f ? _GEN_102 : _GEN_101; // @[lut_mem_online.scala 235:34]
  wire  _GEN_104 = ~io_inputBit ? 1'h0 : _GEN_103; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_105 = _GEN_6084 == 9'h10c ? _GEN_104 : _GEN_103; // @[lut_mem_online.scala 235:34]
  wire  _GEN_106 = ~io_inputBit | _GEN_105; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_107 = _GEN_6084 == 9'h110 ? _GEN_106 : _GEN_105; // @[lut_mem_online.scala 235:34]
  wire  _GEN_108 = ~io_inputBit ? 1'h0 : _GEN_107; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_109 = _GEN_6084 == 9'h114 ? _GEN_108 : _GEN_107; // @[lut_mem_online.scala 235:34]
  wire  _GEN_110 = ~io_inputBit | _GEN_109; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_111 = _GEN_6084 == 9'h118 ? _GEN_110 : _GEN_109; // @[lut_mem_online.scala 235:34]
  wire  _GEN_112 = ~io_inputBit ? 1'h0 : _GEN_111; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_113 = _GEN_6084 == 9'h11c ? _GEN_112 : _GEN_111; // @[lut_mem_online.scala 235:34]
  wire  _GEN_114 = ~io_inputBit | _GEN_113; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_115 = _GEN_6084 == 9'h120 ? _GEN_114 : _GEN_113; // @[lut_mem_online.scala 235:34]
  wire  _GEN_116 = ~io_inputBit ? 1'h0 : _GEN_115; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_117 = _GEN_6085 == 10'h21a ? _GEN_116 : _GEN_115; // @[lut_mem_online.scala 235:34]
  wire  _GEN_118 = io_inputBit | _GEN_117; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_119 = _GEN_6085 == 10'h21a ? _GEN_118 : _GEN_117; // @[lut_mem_online.scala 235:34]
  wire  _GEN_120 = ~io_inputBit | _GEN_119; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_121 = _GEN_6085 == 10'h222 ? _GEN_120 : _GEN_119; // @[lut_mem_online.scala 235:34]
  wire  _GEN_122 = io_inputBit ? 1'h0 : _GEN_121; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_123 = _GEN_6085 == 10'h222 ? _GEN_122 : _GEN_121; // @[lut_mem_online.scala 235:34]
  wire  _GEN_124 = ~io_inputBit ? 1'h0 : _GEN_123; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_125 = _GEN_6085 == 10'h22a ? _GEN_124 : _GEN_123; // @[lut_mem_online.scala 235:34]
  wire  _GEN_126 = io_inputBit | _GEN_125; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_127 = _GEN_6085 == 10'h22a ? _GEN_126 : _GEN_125; // @[lut_mem_online.scala 235:34]
  wire  _GEN_128 = ~io_inputBit | _GEN_127; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_129 = _GEN_6085 == 10'h232 ? _GEN_128 : _GEN_127; // @[lut_mem_online.scala 235:34]
  wire  _GEN_130 = io_inputBit ? 1'h0 : _GEN_129; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_131 = _GEN_6085 == 10'h232 ? _GEN_130 : _GEN_129; // @[lut_mem_online.scala 235:34]
  wire  _GEN_132 = ~io_inputBit ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_133 = _GEN_6085 == 10'h23a ? _GEN_132 : _GEN_131; // @[lut_mem_online.scala 235:34]
  wire  _GEN_134 = io_inputBit | _GEN_133; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_135 = _GEN_6085 == 10'h23a ? _GEN_134 : _GEN_133; // @[lut_mem_online.scala 235:34]
  wire  _GEN_136 = ~io_inputBit | _GEN_135; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_137 = _GEN_6085 == 10'h242 ? _GEN_136 : _GEN_135; // @[lut_mem_online.scala 235:34]
  wire  _GEN_138 = io_inputBit ? 1'h0 : _GEN_137; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_139 = _GEN_6085 == 10'h242 ? _GEN_138 : _GEN_137; // @[lut_mem_online.scala 235:34]
  wire  _GEN_140 = io_inputBit ? 1'h0 : buffer_3; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_141 = i == 8'h0 ? _GEN_140 : buffer_3; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_142 = io_inputBit ? 1'h0 : _GEN_141; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_143 = i == 8'h1 ? _GEN_142 : _GEN_141; // @[lut_mem_online.scala 235:34]
  wire  _GEN_144 = io_inputBit ? 1'h0 : _GEN_143; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_145 = i == 8'h8 ? _GEN_144 : _GEN_143; // @[lut_mem_online.scala 235:34]
  wire  _GEN_146 = ~io_inputBit ? 1'h0 : _GEN_145; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_147 = i == 8'hf ? _GEN_146 : _GEN_145; // @[lut_mem_online.scala 235:34]
  wire  _GEN_148 = io_inputBit ? 1'h0 : _GEN_147; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_149 = i == 8'h11 ? _GEN_148 : _GEN_147; // @[lut_mem_online.scala 235:34]
  wire  _GEN_150 = ~io_inputBit ? 1'h0 : _GEN_149; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_151 = i == 8'h20 ? _GEN_150 : _GEN_149; // @[lut_mem_online.scala 235:34]
  wire  _GEN_152 = io_inputBit ? 1'h0 : _GEN_151; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_153 = i == 8'h23 ? _GEN_152 : _GEN_151; // @[lut_mem_online.scala 235:34]
  wire  _GEN_154 = ~io_inputBit ? 1'h0 : _GEN_153; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_155 = i == 8'h85 ? _GEN_154 : _GEN_153; // @[lut_mem_online.scala 235:34]
  wire  _GEN_156 = ~io_inputBit | _GEN_155; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_157 = i == 8'h86 ? _GEN_156 : _GEN_155; // @[lut_mem_online.scala 235:34]
  wire  _GEN_158 = ~io_inputBit ? 1'h0 : _GEN_157; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_159 = i == 8'h87 ? _GEN_158 : _GEN_157; // @[lut_mem_online.scala 235:34]
  wire  _GEN_160 = ~io_inputBit | _GEN_159; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_161 = i == 8'h88 ? _GEN_160 : _GEN_159; // @[lut_mem_online.scala 235:34]
  wire  _GEN_162 = ~io_inputBit ? 1'h0 : _GEN_161; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_163 = i == 8'h89 ? _GEN_162 : _GEN_161; // @[lut_mem_online.scala 235:34]
  wire  _GEN_164 = ~io_inputBit | _GEN_163; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_165 = i == 8'h8a ? _GEN_164 : _GEN_163; // @[lut_mem_online.scala 235:34]
  wire  _GEN_166 = ~io_inputBit ? 1'h0 : _GEN_165; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_167 = i == 8'h8b ? _GEN_166 : _GEN_165; // @[lut_mem_online.scala 235:34]
  wire  _GEN_168 = ~io_inputBit | _GEN_167; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_169 = i == 8'h8c ? _GEN_168 : _GEN_167; // @[lut_mem_online.scala 235:34]
  wire  _GEN_170 = ~io_inputBit ? 1'h0 : _GEN_169; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_171 = i == 8'h8d ? _GEN_170 : _GEN_169; // @[lut_mem_online.scala 235:34]
  wire  _GEN_172 = ~io_inputBit | _GEN_171; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_173 = i == 8'h8e ? _GEN_172 : _GEN_171; // @[lut_mem_online.scala 235:34]
  wire  _GEN_174 = ~io_inputBit ? 1'h0 : _GEN_173; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_175 = i == 8'h8f ? _GEN_174 : _GEN_173; // @[lut_mem_online.scala 235:34]
  wire  _GEN_176 = ~io_inputBit | _GEN_175; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_177 = i == 8'h90 ? _GEN_176 : _GEN_175; // @[lut_mem_online.scala 235:34]
  wire  _GEN_178 = ~io_inputBit ? 1'h0 : _GEN_177; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_179 = _GEN_6084 == 9'h10c ? _GEN_178 : _GEN_177; // @[lut_mem_online.scala 235:34]
  wire  _GEN_180 = ~io_inputBit | _GEN_179; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_181 = _GEN_6084 == 9'h10e ? _GEN_180 : _GEN_179; // @[lut_mem_online.scala 235:34]
  wire  _GEN_182 = ~io_inputBit ? 1'h0 : _GEN_181; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_183 = _GEN_6084 == 9'h110 ? _GEN_182 : _GEN_181; // @[lut_mem_online.scala 235:34]
  wire  _GEN_184 = ~io_inputBit | _GEN_183; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_185 = _GEN_6084 == 9'h112 ? _GEN_184 : _GEN_183; // @[lut_mem_online.scala 235:34]
  wire  _GEN_186 = ~io_inputBit ? 1'h0 : _GEN_185; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_187 = _GEN_6084 == 9'h114 ? _GEN_186 : _GEN_185; // @[lut_mem_online.scala 235:34]
  wire  _GEN_188 = ~io_inputBit | _GEN_187; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_189 = _GEN_6084 == 9'h116 ? _GEN_188 : _GEN_187; // @[lut_mem_online.scala 235:34]
  wire  _GEN_190 = ~io_inputBit ? 1'h0 : _GEN_189; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_191 = _GEN_6084 == 9'h118 ? _GEN_190 : _GEN_189; // @[lut_mem_online.scala 235:34]
  wire  _GEN_192 = ~io_inputBit | _GEN_191; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_193 = _GEN_6084 == 9'h11a ? _GEN_192 : _GEN_191; // @[lut_mem_online.scala 235:34]
  wire  _GEN_194 = ~io_inputBit ? 1'h0 : _GEN_193; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_195 = _GEN_6084 == 9'h11c ? _GEN_194 : _GEN_193; // @[lut_mem_online.scala 235:34]
  wire  _GEN_196 = ~io_inputBit | _GEN_195; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_197 = _GEN_6084 == 9'h11e ? _GEN_196 : _GEN_195; // @[lut_mem_online.scala 235:34]
  wire  _GEN_198 = ~io_inputBit ? 1'h0 : _GEN_197; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_199 = _GEN_6084 == 9'h120 ? _GEN_198 : _GEN_197; // @[lut_mem_online.scala 235:34]
  wire  _GEN_200 = ~io_inputBit | _GEN_199; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_201 = _GEN_6084 == 9'h122 ? _GEN_200 : _GEN_199; // @[lut_mem_online.scala 235:34]
  wire  _GEN_202 = ~io_inputBit ? 1'h0 : _GEN_201; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_203 = _GEN_6085 == 10'h21a ? _GEN_202 : _GEN_201; // @[lut_mem_online.scala 235:34]
  wire  _GEN_204 = io_inputBit | _GEN_203; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_205 = _GEN_6085 == 10'h21a ? _GEN_204 : _GEN_203; // @[lut_mem_online.scala 235:34]
  wire  _GEN_206 = ~io_inputBit | _GEN_205; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_207 = _GEN_6085 == 10'h21e ? _GEN_206 : _GEN_205; // @[lut_mem_online.scala 235:34]
  wire  _GEN_208 = io_inputBit ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_209 = _GEN_6085 == 10'h21e ? _GEN_208 : _GEN_207; // @[lut_mem_online.scala 235:34]
  wire  _GEN_210 = ~io_inputBit ? 1'h0 : _GEN_209; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_211 = _GEN_6085 == 10'h222 ? _GEN_210 : _GEN_209; // @[lut_mem_online.scala 235:34]
  wire  _GEN_212 = io_inputBit | _GEN_211; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_213 = _GEN_6085 == 10'h222 ? _GEN_212 : _GEN_211; // @[lut_mem_online.scala 235:34]
  wire  _GEN_214 = ~io_inputBit | _GEN_213; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_215 = _GEN_6085 == 10'h226 ? _GEN_214 : _GEN_213; // @[lut_mem_online.scala 235:34]
  wire  _GEN_216 = io_inputBit ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_217 = _GEN_6085 == 10'h226 ? _GEN_216 : _GEN_215; // @[lut_mem_online.scala 235:34]
  wire  _GEN_218 = ~io_inputBit ? 1'h0 : _GEN_217; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_219 = _GEN_6085 == 10'h22a ? _GEN_218 : _GEN_217; // @[lut_mem_online.scala 235:34]
  wire  _GEN_220 = io_inputBit | _GEN_219; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_221 = _GEN_6085 == 10'h22a ? _GEN_220 : _GEN_219; // @[lut_mem_online.scala 235:34]
  wire  _GEN_222 = ~io_inputBit | _GEN_221; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_223 = _GEN_6085 == 10'h22e ? _GEN_222 : _GEN_221; // @[lut_mem_online.scala 235:34]
  wire  _GEN_224 = io_inputBit ? 1'h0 : _GEN_223; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_225 = _GEN_6085 == 10'h22e ? _GEN_224 : _GEN_223; // @[lut_mem_online.scala 235:34]
  wire  _GEN_226 = ~io_inputBit ? 1'h0 : _GEN_225; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_227 = _GEN_6085 == 10'h232 ? _GEN_226 : _GEN_225; // @[lut_mem_online.scala 235:34]
  wire  _GEN_228 = io_inputBit | _GEN_227; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_229 = _GEN_6085 == 10'h232 ? _GEN_228 : _GEN_227; // @[lut_mem_online.scala 235:34]
  wire  _GEN_230 = ~io_inputBit | _GEN_229; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_231 = _GEN_6085 == 10'h236 ? _GEN_230 : _GEN_229; // @[lut_mem_online.scala 235:34]
  wire  _GEN_232 = io_inputBit ? 1'h0 : _GEN_231; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_233 = _GEN_6085 == 10'h236 ? _GEN_232 : _GEN_231; // @[lut_mem_online.scala 235:34]
  wire  _GEN_234 = ~io_inputBit ? 1'h0 : _GEN_233; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_235 = _GEN_6085 == 10'h23a ? _GEN_234 : _GEN_233; // @[lut_mem_online.scala 235:34]
  wire  _GEN_236 = io_inputBit | _GEN_235; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_237 = _GEN_6085 == 10'h23a ? _GEN_236 : _GEN_235; // @[lut_mem_online.scala 235:34]
  wire  _GEN_238 = ~io_inputBit | _GEN_237; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_239 = _GEN_6085 == 10'h23e ? _GEN_238 : _GEN_237; // @[lut_mem_online.scala 235:34]
  wire  _GEN_240 = io_inputBit ? 1'h0 : _GEN_239; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_241 = _GEN_6085 == 10'h23e ? _GEN_240 : _GEN_239; // @[lut_mem_online.scala 235:34]
  wire  _GEN_242 = ~io_inputBit ? 1'h0 : _GEN_241; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_243 = _GEN_6085 == 10'h242 ? _GEN_242 : _GEN_241; // @[lut_mem_online.scala 235:34]
  wire  _GEN_244 = io_inputBit | _GEN_243; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_245 = _GEN_6085 == 10'h242 ? _GEN_244 : _GEN_243; // @[lut_mem_online.scala 235:34]
  wire  _GEN_246 = ~io_inputBit | _GEN_245; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_247 = _GEN_6085 == 10'h246 ? _GEN_246 : _GEN_245; // @[lut_mem_online.scala 235:34]
  wire  _GEN_248 = io_inputBit ? 1'h0 : _GEN_247; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_249 = _GEN_6085 == 10'h246 ? _GEN_248 : _GEN_247; // @[lut_mem_online.scala 235:34]
  wire  _GEN_250 = io_inputBit ? 1'h0 : buffer_4; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_251 = i == 8'h0 ? _GEN_250 : buffer_4; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_252 = io_inputBit ? 1'h0 : _GEN_251; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_253 = i == 8'h1 ? _GEN_252 : _GEN_251; // @[lut_mem_online.scala 235:34]
  wire  _GEN_254 = io_inputBit ? 1'h0 : _GEN_253; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_255 = i == 8'h8 ? _GEN_254 : _GEN_253; // @[lut_mem_online.scala 235:34]
  wire  _GEN_256 = ~io_inputBit | _GEN_255; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_257 = i == 8'hf ? _GEN_256 : _GEN_255; // @[lut_mem_online.scala 235:34]
  wire  _GEN_258 = io_inputBit ? 1'h0 : _GEN_257; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_259 = i == 8'h11 ? _GEN_258 : _GEN_257; // @[lut_mem_online.scala 235:34]
  wire  _GEN_260 = ~io_inputBit | _GEN_259; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_261 = i == 8'h20 ? _GEN_260 : _GEN_259; // @[lut_mem_online.scala 235:34]
  wire  _GEN_262 = io_inputBit ? 1'h0 : _GEN_261; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_263 = i == 8'h48 ? _GEN_262 : _GEN_261; // @[lut_mem_online.scala 235:34]
  wire  _GEN_264 = io_inputBit ? 1'h0 : _GEN_263; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_265 = i == 8'h91 ? _GEN_264 : _GEN_263; // @[lut_mem_online.scala 235:34]
  wire  _GEN_266 = ~io_inputBit | _GEN_265; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_267 = _GEN_6084 == 9'h10b ? _GEN_266 : _GEN_265; // @[lut_mem_online.scala 235:34]
  wire  _GEN_268 = ~io_inputBit ? 1'h0 : _GEN_267; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_269 = _GEN_6084 == 9'h10c ? _GEN_268 : _GEN_267; // @[lut_mem_online.scala 235:34]
  wire  _GEN_270 = ~io_inputBit | _GEN_269; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_271 = _GEN_6084 == 9'h10d ? _GEN_270 : _GEN_269; // @[lut_mem_online.scala 235:34]
  wire  _GEN_272 = ~io_inputBit ? 1'h0 : _GEN_271; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_273 = _GEN_6084 == 9'h10e ? _GEN_272 : _GEN_271; // @[lut_mem_online.scala 235:34]
  wire  _GEN_274 = ~io_inputBit | _GEN_273; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_275 = _GEN_6084 == 9'h10f ? _GEN_274 : _GEN_273; // @[lut_mem_online.scala 235:34]
  wire  _GEN_276 = ~io_inputBit ? 1'h0 : _GEN_275; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_277 = _GEN_6084 == 9'h110 ? _GEN_276 : _GEN_275; // @[lut_mem_online.scala 235:34]
  wire  _GEN_278 = ~io_inputBit | _GEN_277; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_279 = _GEN_6084 == 9'h111 ? _GEN_278 : _GEN_277; // @[lut_mem_online.scala 235:34]
  wire  _GEN_280 = ~io_inputBit ? 1'h0 : _GEN_279; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_281 = _GEN_6084 == 9'h112 ? _GEN_280 : _GEN_279; // @[lut_mem_online.scala 235:34]
  wire  _GEN_282 = ~io_inputBit | _GEN_281; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_283 = _GEN_6084 == 9'h113 ? _GEN_282 : _GEN_281; // @[lut_mem_online.scala 235:34]
  wire  _GEN_284 = ~io_inputBit ? 1'h0 : _GEN_283; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_285 = _GEN_6084 == 9'h114 ? _GEN_284 : _GEN_283; // @[lut_mem_online.scala 235:34]
  wire  _GEN_286 = ~io_inputBit | _GEN_285; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_287 = _GEN_6084 == 9'h115 ? _GEN_286 : _GEN_285; // @[lut_mem_online.scala 235:34]
  wire  _GEN_288 = ~io_inputBit ? 1'h0 : _GEN_287; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_289 = _GEN_6084 == 9'h116 ? _GEN_288 : _GEN_287; // @[lut_mem_online.scala 235:34]
  wire  _GEN_290 = ~io_inputBit | _GEN_289; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_291 = _GEN_6084 == 9'h117 ? _GEN_290 : _GEN_289; // @[lut_mem_online.scala 235:34]
  wire  _GEN_292 = ~io_inputBit ? 1'h0 : _GEN_291; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_293 = _GEN_6084 == 9'h118 ? _GEN_292 : _GEN_291; // @[lut_mem_online.scala 235:34]
  wire  _GEN_294 = ~io_inputBit | _GEN_293; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_295 = _GEN_6084 == 9'h119 ? _GEN_294 : _GEN_293; // @[lut_mem_online.scala 235:34]
  wire  _GEN_296 = ~io_inputBit ? 1'h0 : _GEN_295; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_297 = _GEN_6084 == 9'h11a ? _GEN_296 : _GEN_295; // @[lut_mem_online.scala 235:34]
  wire  _GEN_298 = ~io_inputBit | _GEN_297; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_299 = _GEN_6084 == 9'h11b ? _GEN_298 : _GEN_297; // @[lut_mem_online.scala 235:34]
  wire  _GEN_300 = ~io_inputBit ? 1'h0 : _GEN_299; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_301 = _GEN_6084 == 9'h11c ? _GEN_300 : _GEN_299; // @[lut_mem_online.scala 235:34]
  wire  _GEN_302 = ~io_inputBit | _GEN_301; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_303 = _GEN_6084 == 9'h11d ? _GEN_302 : _GEN_301; // @[lut_mem_online.scala 235:34]
  wire  _GEN_304 = ~io_inputBit ? 1'h0 : _GEN_303; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_305 = _GEN_6084 == 9'h11e ? _GEN_304 : _GEN_303; // @[lut_mem_online.scala 235:34]
  wire  _GEN_306 = ~io_inputBit | _GEN_305; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_307 = _GEN_6084 == 9'h11f ? _GEN_306 : _GEN_305; // @[lut_mem_online.scala 235:34]
  wire  _GEN_308 = ~io_inputBit ? 1'h0 : _GEN_307; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_309 = _GEN_6084 == 9'h120 ? _GEN_308 : _GEN_307; // @[lut_mem_online.scala 235:34]
  wire  _GEN_310 = ~io_inputBit | _GEN_309; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_311 = _GEN_6084 == 9'h121 ? _GEN_310 : _GEN_309; // @[lut_mem_online.scala 235:34]
  wire  _GEN_312 = ~io_inputBit ? 1'h0 : _GEN_311; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_313 = _GEN_6084 == 9'h122 ? _GEN_312 : _GEN_311; // @[lut_mem_online.scala 235:34]
  wire  _GEN_314 = ~io_inputBit | _GEN_313; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_315 = _GEN_6084 == 9'h123 ? _GEN_314 : _GEN_313; // @[lut_mem_online.scala 235:34]
  wire  _GEN_316 = ~io_inputBit | _GEN_315; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_317 = _GEN_6085 == 10'h218 ? _GEN_316 : _GEN_315; // @[lut_mem_online.scala 235:34]
  wire  _GEN_318 = io_inputBit ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_319 = _GEN_6085 == 10'h218 ? _GEN_318 : _GEN_317; // @[lut_mem_online.scala 235:34]
  wire  _GEN_320 = ~io_inputBit ? 1'h0 : _GEN_319; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_321 = _GEN_6085 == 10'h21a ? _GEN_320 : _GEN_319; // @[lut_mem_online.scala 235:34]
  wire  _GEN_322 = io_inputBit | _GEN_321; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_323 = _GEN_6085 == 10'h21a ? _GEN_322 : _GEN_321; // @[lut_mem_online.scala 235:34]
  wire  _GEN_324 = ~io_inputBit | _GEN_323; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_325 = _GEN_6085 == 10'h21c ? _GEN_324 : _GEN_323; // @[lut_mem_online.scala 235:34]
  wire  _GEN_326 = io_inputBit ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_327 = _GEN_6085 == 10'h21c ? _GEN_326 : _GEN_325; // @[lut_mem_online.scala 235:34]
  wire  _GEN_328 = ~io_inputBit ? 1'h0 : _GEN_327; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_329 = _GEN_6085 == 10'h21e ? _GEN_328 : _GEN_327; // @[lut_mem_online.scala 235:34]
  wire  _GEN_330 = io_inputBit | _GEN_329; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_331 = _GEN_6085 == 10'h21e ? _GEN_330 : _GEN_329; // @[lut_mem_online.scala 235:34]
  wire  _GEN_332 = ~io_inputBit | _GEN_331; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_333 = _GEN_6085 == 10'h220 ? _GEN_332 : _GEN_331; // @[lut_mem_online.scala 235:34]
  wire  _GEN_334 = io_inputBit ? 1'h0 : _GEN_333; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_335 = _GEN_6085 == 10'h220 ? _GEN_334 : _GEN_333; // @[lut_mem_online.scala 235:34]
  wire  _GEN_336 = ~io_inputBit ? 1'h0 : _GEN_335; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_337 = _GEN_6085 == 10'h222 ? _GEN_336 : _GEN_335; // @[lut_mem_online.scala 235:34]
  wire  _GEN_338 = io_inputBit | _GEN_337; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_339 = _GEN_6085 == 10'h222 ? _GEN_338 : _GEN_337; // @[lut_mem_online.scala 235:34]
  wire  _GEN_340 = ~io_inputBit | _GEN_339; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_341 = _GEN_6085 == 10'h224 ? _GEN_340 : _GEN_339; // @[lut_mem_online.scala 235:34]
  wire  _GEN_342 = io_inputBit ? 1'h0 : _GEN_341; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_343 = _GEN_6085 == 10'h224 ? _GEN_342 : _GEN_341; // @[lut_mem_online.scala 235:34]
  wire  _GEN_344 = ~io_inputBit ? 1'h0 : _GEN_343; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_345 = _GEN_6085 == 10'h226 ? _GEN_344 : _GEN_343; // @[lut_mem_online.scala 235:34]
  wire  _GEN_346 = io_inputBit | _GEN_345; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_347 = _GEN_6085 == 10'h226 ? _GEN_346 : _GEN_345; // @[lut_mem_online.scala 235:34]
  wire  _GEN_348 = ~io_inputBit | _GEN_347; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_349 = _GEN_6085 == 10'h228 ? _GEN_348 : _GEN_347; // @[lut_mem_online.scala 235:34]
  wire  _GEN_350 = io_inputBit ? 1'h0 : _GEN_349; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_351 = _GEN_6085 == 10'h228 ? _GEN_350 : _GEN_349; // @[lut_mem_online.scala 235:34]
  wire  _GEN_352 = ~io_inputBit ? 1'h0 : _GEN_351; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_353 = _GEN_6085 == 10'h22a ? _GEN_352 : _GEN_351; // @[lut_mem_online.scala 235:34]
  wire  _GEN_354 = io_inputBit | _GEN_353; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_355 = _GEN_6085 == 10'h22a ? _GEN_354 : _GEN_353; // @[lut_mem_online.scala 235:34]
  wire  _GEN_356 = ~io_inputBit | _GEN_355; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_357 = _GEN_6085 == 10'h22c ? _GEN_356 : _GEN_355; // @[lut_mem_online.scala 235:34]
  wire  _GEN_358 = io_inputBit ? 1'h0 : _GEN_357; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_359 = _GEN_6085 == 10'h22c ? _GEN_358 : _GEN_357; // @[lut_mem_online.scala 235:34]
  wire  _GEN_360 = ~io_inputBit ? 1'h0 : _GEN_359; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_361 = _GEN_6085 == 10'h22e ? _GEN_360 : _GEN_359; // @[lut_mem_online.scala 235:34]
  wire  _GEN_362 = io_inputBit | _GEN_361; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_363 = _GEN_6085 == 10'h22e ? _GEN_362 : _GEN_361; // @[lut_mem_online.scala 235:34]
  wire  _GEN_364 = ~io_inputBit | _GEN_363; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_365 = _GEN_6085 == 10'h230 ? _GEN_364 : _GEN_363; // @[lut_mem_online.scala 235:34]
  wire  _GEN_366 = io_inputBit ? 1'h0 : _GEN_365; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_367 = _GEN_6085 == 10'h230 ? _GEN_366 : _GEN_365; // @[lut_mem_online.scala 235:34]
  wire  _GEN_368 = ~io_inputBit ? 1'h0 : _GEN_367; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_369 = _GEN_6085 == 10'h232 ? _GEN_368 : _GEN_367; // @[lut_mem_online.scala 235:34]
  wire  _GEN_370 = io_inputBit | _GEN_369; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_371 = _GEN_6085 == 10'h232 ? _GEN_370 : _GEN_369; // @[lut_mem_online.scala 235:34]
  wire  _GEN_372 = ~io_inputBit | _GEN_371; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_373 = _GEN_6085 == 10'h234 ? _GEN_372 : _GEN_371; // @[lut_mem_online.scala 235:34]
  wire  _GEN_374 = io_inputBit ? 1'h0 : _GEN_373; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_375 = _GEN_6085 == 10'h234 ? _GEN_374 : _GEN_373; // @[lut_mem_online.scala 235:34]
  wire  _GEN_376 = ~io_inputBit ? 1'h0 : _GEN_375; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_377 = _GEN_6085 == 10'h236 ? _GEN_376 : _GEN_375; // @[lut_mem_online.scala 235:34]
  wire  _GEN_378 = io_inputBit | _GEN_377; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_379 = _GEN_6085 == 10'h236 ? _GEN_378 : _GEN_377; // @[lut_mem_online.scala 235:34]
  wire  _GEN_380 = ~io_inputBit | _GEN_379; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_381 = _GEN_6085 == 10'h238 ? _GEN_380 : _GEN_379; // @[lut_mem_online.scala 235:34]
  wire  _GEN_382 = io_inputBit ? 1'h0 : _GEN_381; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_383 = _GEN_6085 == 10'h238 ? _GEN_382 : _GEN_381; // @[lut_mem_online.scala 235:34]
  wire  _GEN_384 = ~io_inputBit ? 1'h0 : _GEN_383; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_385 = _GEN_6085 == 10'h23a ? _GEN_384 : _GEN_383; // @[lut_mem_online.scala 235:34]
  wire  _GEN_386 = io_inputBit | _GEN_385; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_387 = _GEN_6085 == 10'h23a ? _GEN_386 : _GEN_385; // @[lut_mem_online.scala 235:34]
  wire  _GEN_388 = ~io_inputBit | _GEN_387; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_389 = _GEN_6085 == 10'h23c ? _GEN_388 : _GEN_387; // @[lut_mem_online.scala 235:34]
  wire  _GEN_390 = io_inputBit ? 1'h0 : _GEN_389; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_391 = _GEN_6085 == 10'h23c ? _GEN_390 : _GEN_389; // @[lut_mem_online.scala 235:34]
  wire  _GEN_392 = ~io_inputBit ? 1'h0 : _GEN_391; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_393 = _GEN_6085 == 10'h23e ? _GEN_392 : _GEN_391; // @[lut_mem_online.scala 235:34]
  wire  _GEN_394 = io_inputBit | _GEN_393; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_395 = _GEN_6085 == 10'h23e ? _GEN_394 : _GEN_393; // @[lut_mem_online.scala 235:34]
  wire  _GEN_396 = ~io_inputBit | _GEN_395; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_397 = _GEN_6085 == 10'h240 ? _GEN_396 : _GEN_395; // @[lut_mem_online.scala 235:34]
  wire  _GEN_398 = io_inputBit ? 1'h0 : _GEN_397; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_399 = _GEN_6085 == 10'h240 ? _GEN_398 : _GEN_397; // @[lut_mem_online.scala 235:34]
  wire  _GEN_400 = ~io_inputBit ? 1'h0 : _GEN_399; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_401 = _GEN_6085 == 10'h242 ? _GEN_400 : _GEN_399; // @[lut_mem_online.scala 235:34]
  wire  _GEN_402 = io_inputBit | _GEN_401; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_403 = _GEN_6085 == 10'h242 ? _GEN_402 : _GEN_401; // @[lut_mem_online.scala 235:34]
  wire  _GEN_404 = ~io_inputBit | _GEN_403; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_405 = _GEN_6085 == 10'h244 ? _GEN_404 : _GEN_403; // @[lut_mem_online.scala 235:34]
  wire  _GEN_406 = io_inputBit ? 1'h0 : _GEN_405; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_407 = _GEN_6085 == 10'h244 ? _GEN_406 : _GEN_405; // @[lut_mem_online.scala 235:34]
  wire  _GEN_408 = ~io_inputBit ? 1'h0 : _GEN_407; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_409 = _GEN_6085 == 10'h246 ? _GEN_408 : _GEN_407; // @[lut_mem_online.scala 235:34]
  wire  _GEN_410 = io_inputBit | _GEN_409; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_411 = _GEN_6085 == 10'h246 ? _GEN_410 : _GEN_409; // @[lut_mem_online.scala 235:34]
  wire  _GEN_412 = ~io_inputBit | _GEN_411; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_413 = _GEN_6085 == 10'h248 ? _GEN_412 : _GEN_411; // @[lut_mem_online.scala 235:34]
  wire  _GEN_414 = io_inputBit ? 1'h0 : _GEN_413; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_415 = _GEN_6085 == 10'h248 ? _GEN_414 : _GEN_413; // @[lut_mem_online.scala 235:34]
  wire  _GEN_416 = io_inputBit ? 1'h0 : buffer_5; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_417 = i == 8'h0 ? _GEN_416 : buffer_5; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_418 = io_inputBit ? 1'h0 : _GEN_417; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_419 = i == 8'h1 ? _GEN_418 : _GEN_417; // @[lut_mem_online.scala 235:34]
  wire  _GEN_420 = io_inputBit ? 1'h0 : _GEN_419; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_421 = i == 8'h8 ? _GEN_420 : _GEN_419; // @[lut_mem_online.scala 235:34]
  wire  _GEN_422 = ~io_inputBit ? 1'h0 : _GEN_421; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_423 = i == 8'hf ? _GEN_422 : _GEN_421; // @[lut_mem_online.scala 235:34]
  wire  _GEN_424 = io_inputBit ? 1'h0 : _GEN_423; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_425 = i == 8'h11 ? _GEN_424 : _GEN_423; // @[lut_mem_online.scala 235:34]
  wire  _GEN_426 = ~io_inputBit ? 1'h0 : _GEN_425; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_427 = i == 8'h20 ? _GEN_426 : _GEN_425; // @[lut_mem_online.scala 235:34]
  wire  _GEN_428 = io_inputBit ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_429 = i == 8'h48 ? _GEN_428 : _GEN_427; // @[lut_mem_online.scala 235:34]
  wire  _GEN_430 = ~io_inputBit ? 1'h0 : _GEN_429; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_431 = _GEN_6084 == 9'h10b ? _GEN_430 : _GEN_429; // @[lut_mem_online.scala 235:34]
  wire  _GEN_432 = io_inputBit ? 1'h0 : _GEN_431; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_433 = _GEN_6084 == 9'h124 ? _GEN_432 : _GEN_431; // @[lut_mem_online.scala 235:34]
  wire  _GEN_434 = ~io_inputBit ? 1'h0 : _GEN_433; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_435 = _GEN_6085 == 10'h218 ? _GEN_434 : _GEN_433; // @[lut_mem_online.scala 235:34]
  wire  _GEN_436 = io_inputBit | _GEN_435; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_437 = _GEN_6085 == 10'h218 ? _GEN_436 : _GEN_435; // @[lut_mem_online.scala 235:34]
  wire  _GEN_438 = ~io_inputBit | _GEN_437; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_439 = _GEN_6085 == 10'h219 ? _GEN_438 : _GEN_437; // @[lut_mem_online.scala 235:34]
  wire  _GEN_440 = io_inputBit ? 1'h0 : _GEN_439; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_441 = _GEN_6085 == 10'h219 ? _GEN_440 : _GEN_439; // @[lut_mem_online.scala 235:34]
  wire  _GEN_442 = ~io_inputBit ? 1'h0 : _GEN_441; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_443 = _GEN_6085 == 10'h21a ? _GEN_442 : _GEN_441; // @[lut_mem_online.scala 235:34]
  wire  _GEN_444 = io_inputBit | _GEN_443; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_445 = _GEN_6085 == 10'h21a ? _GEN_444 : _GEN_443; // @[lut_mem_online.scala 235:34]
  wire  _GEN_446 = ~io_inputBit | _GEN_445; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_447 = _GEN_6085 == 10'h21b ? _GEN_446 : _GEN_445; // @[lut_mem_online.scala 235:34]
  wire  _GEN_448 = io_inputBit ? 1'h0 : _GEN_447; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_449 = _GEN_6085 == 10'h21b ? _GEN_448 : _GEN_447; // @[lut_mem_online.scala 235:34]
  wire  _GEN_450 = ~io_inputBit ? 1'h0 : _GEN_449; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_451 = _GEN_6085 == 10'h21c ? _GEN_450 : _GEN_449; // @[lut_mem_online.scala 235:34]
  wire  _GEN_452 = io_inputBit | _GEN_451; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_453 = _GEN_6085 == 10'h21c ? _GEN_452 : _GEN_451; // @[lut_mem_online.scala 235:34]
  wire  _GEN_454 = ~io_inputBit | _GEN_453; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_455 = _GEN_6085 == 10'h21d ? _GEN_454 : _GEN_453; // @[lut_mem_online.scala 235:34]
  wire  _GEN_456 = io_inputBit ? 1'h0 : _GEN_455; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_457 = _GEN_6085 == 10'h21d ? _GEN_456 : _GEN_455; // @[lut_mem_online.scala 235:34]
  wire  _GEN_458 = ~io_inputBit ? 1'h0 : _GEN_457; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_459 = _GEN_6085 == 10'h21e ? _GEN_458 : _GEN_457; // @[lut_mem_online.scala 235:34]
  wire  _GEN_460 = io_inputBit | _GEN_459; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_461 = _GEN_6085 == 10'h21e ? _GEN_460 : _GEN_459; // @[lut_mem_online.scala 235:34]
  wire  _GEN_462 = ~io_inputBit | _GEN_461; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_463 = _GEN_6085 == 10'h21f ? _GEN_462 : _GEN_461; // @[lut_mem_online.scala 235:34]
  wire  _GEN_464 = io_inputBit ? 1'h0 : _GEN_463; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_465 = _GEN_6085 == 10'h21f ? _GEN_464 : _GEN_463; // @[lut_mem_online.scala 235:34]
  wire  _GEN_466 = ~io_inputBit ? 1'h0 : _GEN_465; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_467 = _GEN_6085 == 10'h220 ? _GEN_466 : _GEN_465; // @[lut_mem_online.scala 235:34]
  wire  _GEN_468 = io_inputBit | _GEN_467; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_469 = _GEN_6085 == 10'h220 ? _GEN_468 : _GEN_467; // @[lut_mem_online.scala 235:34]
  wire  _GEN_470 = ~io_inputBit | _GEN_469; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_471 = _GEN_6085 == 10'h221 ? _GEN_470 : _GEN_469; // @[lut_mem_online.scala 235:34]
  wire  _GEN_472 = io_inputBit ? 1'h0 : _GEN_471; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_473 = _GEN_6085 == 10'h221 ? _GEN_472 : _GEN_471; // @[lut_mem_online.scala 235:34]
  wire  _GEN_474 = ~io_inputBit ? 1'h0 : _GEN_473; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_475 = _GEN_6085 == 10'h222 ? _GEN_474 : _GEN_473; // @[lut_mem_online.scala 235:34]
  wire  _GEN_476 = io_inputBit | _GEN_475; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_477 = _GEN_6085 == 10'h222 ? _GEN_476 : _GEN_475; // @[lut_mem_online.scala 235:34]
  wire  _GEN_478 = ~io_inputBit | _GEN_477; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_479 = _GEN_6085 == 10'h223 ? _GEN_478 : _GEN_477; // @[lut_mem_online.scala 235:34]
  wire  _GEN_480 = io_inputBit ? 1'h0 : _GEN_479; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_481 = _GEN_6085 == 10'h223 ? _GEN_480 : _GEN_479; // @[lut_mem_online.scala 235:34]
  wire  _GEN_482 = ~io_inputBit ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_483 = _GEN_6085 == 10'h224 ? _GEN_482 : _GEN_481; // @[lut_mem_online.scala 235:34]
  wire  _GEN_484 = io_inputBit | _GEN_483; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_485 = _GEN_6085 == 10'h224 ? _GEN_484 : _GEN_483; // @[lut_mem_online.scala 235:34]
  wire  _GEN_486 = ~io_inputBit | _GEN_485; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_487 = _GEN_6085 == 10'h225 ? _GEN_486 : _GEN_485; // @[lut_mem_online.scala 235:34]
  wire  _GEN_488 = io_inputBit ? 1'h0 : _GEN_487; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_489 = _GEN_6085 == 10'h225 ? _GEN_488 : _GEN_487; // @[lut_mem_online.scala 235:34]
  wire  _GEN_490 = ~io_inputBit ? 1'h0 : _GEN_489; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_491 = _GEN_6085 == 10'h226 ? _GEN_490 : _GEN_489; // @[lut_mem_online.scala 235:34]
  wire  _GEN_492 = io_inputBit | _GEN_491; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_493 = _GEN_6085 == 10'h226 ? _GEN_492 : _GEN_491; // @[lut_mem_online.scala 235:34]
  wire  _GEN_494 = ~io_inputBit | _GEN_493; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_495 = _GEN_6085 == 10'h227 ? _GEN_494 : _GEN_493; // @[lut_mem_online.scala 235:34]
  wire  _GEN_496 = io_inputBit ? 1'h0 : _GEN_495; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_497 = _GEN_6085 == 10'h227 ? _GEN_496 : _GEN_495; // @[lut_mem_online.scala 235:34]
  wire  _GEN_498 = ~io_inputBit ? 1'h0 : _GEN_497; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_499 = _GEN_6085 == 10'h228 ? _GEN_498 : _GEN_497; // @[lut_mem_online.scala 235:34]
  wire  _GEN_500 = io_inputBit | _GEN_499; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_501 = _GEN_6085 == 10'h228 ? _GEN_500 : _GEN_499; // @[lut_mem_online.scala 235:34]
  wire  _GEN_502 = ~io_inputBit | _GEN_501; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_503 = _GEN_6085 == 10'h229 ? _GEN_502 : _GEN_501; // @[lut_mem_online.scala 235:34]
  wire  _GEN_504 = io_inputBit ? 1'h0 : _GEN_503; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_505 = _GEN_6085 == 10'h229 ? _GEN_504 : _GEN_503; // @[lut_mem_online.scala 235:34]
  wire  _GEN_506 = ~io_inputBit ? 1'h0 : _GEN_505; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_507 = _GEN_6085 == 10'h22a ? _GEN_506 : _GEN_505; // @[lut_mem_online.scala 235:34]
  wire  _GEN_508 = io_inputBit | _GEN_507; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_509 = _GEN_6085 == 10'h22a ? _GEN_508 : _GEN_507; // @[lut_mem_online.scala 235:34]
  wire  _GEN_510 = ~io_inputBit | _GEN_509; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_511 = _GEN_6085 == 10'h22b ? _GEN_510 : _GEN_509; // @[lut_mem_online.scala 235:34]
  wire  _GEN_512 = io_inputBit ? 1'h0 : _GEN_511; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_513 = _GEN_6085 == 10'h22b ? _GEN_512 : _GEN_511; // @[lut_mem_online.scala 235:34]
  wire  _GEN_514 = ~io_inputBit ? 1'h0 : _GEN_513; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_515 = _GEN_6085 == 10'h22c ? _GEN_514 : _GEN_513; // @[lut_mem_online.scala 235:34]
  wire  _GEN_516 = io_inputBit | _GEN_515; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_517 = _GEN_6085 == 10'h22c ? _GEN_516 : _GEN_515; // @[lut_mem_online.scala 235:34]
  wire  _GEN_518 = ~io_inputBit | _GEN_517; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_519 = _GEN_6085 == 10'h22d ? _GEN_518 : _GEN_517; // @[lut_mem_online.scala 235:34]
  wire  _GEN_520 = io_inputBit ? 1'h0 : _GEN_519; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_521 = _GEN_6085 == 10'h22d ? _GEN_520 : _GEN_519; // @[lut_mem_online.scala 235:34]
  wire  _GEN_522 = ~io_inputBit ? 1'h0 : _GEN_521; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_523 = _GEN_6085 == 10'h22e ? _GEN_522 : _GEN_521; // @[lut_mem_online.scala 235:34]
  wire  _GEN_524 = io_inputBit | _GEN_523; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_525 = _GEN_6085 == 10'h22e ? _GEN_524 : _GEN_523; // @[lut_mem_online.scala 235:34]
  wire  _GEN_526 = ~io_inputBit | _GEN_525; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_527 = _GEN_6085 == 10'h22f ? _GEN_526 : _GEN_525; // @[lut_mem_online.scala 235:34]
  wire  _GEN_528 = io_inputBit ? 1'h0 : _GEN_527; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_529 = _GEN_6085 == 10'h22f ? _GEN_528 : _GEN_527; // @[lut_mem_online.scala 235:34]
  wire  _GEN_530 = ~io_inputBit ? 1'h0 : _GEN_529; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_531 = _GEN_6085 == 10'h230 ? _GEN_530 : _GEN_529; // @[lut_mem_online.scala 235:34]
  wire  _GEN_532 = io_inputBit | _GEN_531; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_533 = _GEN_6085 == 10'h230 ? _GEN_532 : _GEN_531; // @[lut_mem_online.scala 235:34]
  wire  _GEN_534 = ~io_inputBit | _GEN_533; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_535 = _GEN_6085 == 10'h231 ? _GEN_534 : _GEN_533; // @[lut_mem_online.scala 235:34]
  wire  _GEN_536 = io_inputBit ? 1'h0 : _GEN_535; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_537 = _GEN_6085 == 10'h231 ? _GEN_536 : _GEN_535; // @[lut_mem_online.scala 235:34]
  wire  _GEN_538 = ~io_inputBit ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_539 = _GEN_6085 == 10'h232 ? _GEN_538 : _GEN_537; // @[lut_mem_online.scala 235:34]
  wire  _GEN_540 = io_inputBit | _GEN_539; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_541 = _GEN_6085 == 10'h232 ? _GEN_540 : _GEN_539; // @[lut_mem_online.scala 235:34]
  wire  _GEN_542 = ~io_inputBit | _GEN_541; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_543 = _GEN_6085 == 10'h233 ? _GEN_542 : _GEN_541; // @[lut_mem_online.scala 235:34]
  wire  _GEN_544 = io_inputBit ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_545 = _GEN_6085 == 10'h233 ? _GEN_544 : _GEN_543; // @[lut_mem_online.scala 235:34]
  wire  _GEN_546 = ~io_inputBit ? 1'h0 : _GEN_545; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_547 = _GEN_6085 == 10'h234 ? _GEN_546 : _GEN_545; // @[lut_mem_online.scala 235:34]
  wire  _GEN_548 = io_inputBit | _GEN_547; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_549 = _GEN_6085 == 10'h234 ? _GEN_548 : _GEN_547; // @[lut_mem_online.scala 235:34]
  wire  _GEN_550 = ~io_inputBit | _GEN_549; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_551 = _GEN_6085 == 10'h235 ? _GEN_550 : _GEN_549; // @[lut_mem_online.scala 235:34]
  wire  _GEN_552 = io_inputBit ? 1'h0 : _GEN_551; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_553 = _GEN_6085 == 10'h235 ? _GEN_552 : _GEN_551; // @[lut_mem_online.scala 235:34]
  wire  _GEN_554 = ~io_inputBit ? 1'h0 : _GEN_553; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_555 = _GEN_6085 == 10'h236 ? _GEN_554 : _GEN_553; // @[lut_mem_online.scala 235:34]
  wire  _GEN_556 = io_inputBit | _GEN_555; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_557 = _GEN_6085 == 10'h236 ? _GEN_556 : _GEN_555; // @[lut_mem_online.scala 235:34]
  wire  _GEN_558 = ~io_inputBit | _GEN_557; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_559 = _GEN_6085 == 10'h237 ? _GEN_558 : _GEN_557; // @[lut_mem_online.scala 235:34]
  wire  _GEN_560 = io_inputBit ? 1'h0 : _GEN_559; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_561 = _GEN_6085 == 10'h237 ? _GEN_560 : _GEN_559; // @[lut_mem_online.scala 235:34]
  wire  _GEN_562 = ~io_inputBit ? 1'h0 : _GEN_561; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_563 = _GEN_6085 == 10'h238 ? _GEN_562 : _GEN_561; // @[lut_mem_online.scala 235:34]
  wire  _GEN_564 = io_inputBit | _GEN_563; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_565 = _GEN_6085 == 10'h238 ? _GEN_564 : _GEN_563; // @[lut_mem_online.scala 235:34]
  wire  _GEN_566 = ~io_inputBit | _GEN_565; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_567 = _GEN_6085 == 10'h239 ? _GEN_566 : _GEN_565; // @[lut_mem_online.scala 235:34]
  wire  _GEN_568 = io_inputBit ? 1'h0 : _GEN_567; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_569 = _GEN_6085 == 10'h239 ? _GEN_568 : _GEN_567; // @[lut_mem_online.scala 235:34]
  wire  _GEN_570 = ~io_inputBit ? 1'h0 : _GEN_569; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_571 = _GEN_6085 == 10'h23a ? _GEN_570 : _GEN_569; // @[lut_mem_online.scala 235:34]
  wire  _GEN_572 = io_inputBit | _GEN_571; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_573 = _GEN_6085 == 10'h23a ? _GEN_572 : _GEN_571; // @[lut_mem_online.scala 235:34]
  wire  _GEN_574 = ~io_inputBit | _GEN_573; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_575 = _GEN_6085 == 10'h23b ? _GEN_574 : _GEN_573; // @[lut_mem_online.scala 235:34]
  wire  _GEN_576 = io_inputBit ? 1'h0 : _GEN_575; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_577 = _GEN_6085 == 10'h23b ? _GEN_576 : _GEN_575; // @[lut_mem_online.scala 235:34]
  wire  _GEN_578 = ~io_inputBit ? 1'h0 : _GEN_577; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_579 = _GEN_6085 == 10'h23c ? _GEN_578 : _GEN_577; // @[lut_mem_online.scala 235:34]
  wire  _GEN_580 = io_inputBit | _GEN_579; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_581 = _GEN_6085 == 10'h23c ? _GEN_580 : _GEN_579; // @[lut_mem_online.scala 235:34]
  wire  _GEN_582 = ~io_inputBit | _GEN_581; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_583 = _GEN_6085 == 10'h23d ? _GEN_582 : _GEN_581; // @[lut_mem_online.scala 235:34]
  wire  _GEN_584 = io_inputBit ? 1'h0 : _GEN_583; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_585 = _GEN_6085 == 10'h23d ? _GEN_584 : _GEN_583; // @[lut_mem_online.scala 235:34]
  wire  _GEN_586 = ~io_inputBit ? 1'h0 : _GEN_585; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_587 = _GEN_6085 == 10'h23e ? _GEN_586 : _GEN_585; // @[lut_mem_online.scala 235:34]
  wire  _GEN_588 = io_inputBit | _GEN_587; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_589 = _GEN_6085 == 10'h23e ? _GEN_588 : _GEN_587; // @[lut_mem_online.scala 235:34]
  wire  _GEN_590 = ~io_inputBit | _GEN_589; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_591 = _GEN_6085 == 10'h23f ? _GEN_590 : _GEN_589; // @[lut_mem_online.scala 235:34]
  wire  _GEN_592 = io_inputBit ? 1'h0 : _GEN_591; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_593 = _GEN_6085 == 10'h23f ? _GEN_592 : _GEN_591; // @[lut_mem_online.scala 235:34]
  wire  _GEN_594 = ~io_inputBit ? 1'h0 : _GEN_593; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_595 = _GEN_6085 == 10'h240 ? _GEN_594 : _GEN_593; // @[lut_mem_online.scala 235:34]
  wire  _GEN_596 = io_inputBit | _GEN_595; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_597 = _GEN_6085 == 10'h240 ? _GEN_596 : _GEN_595; // @[lut_mem_online.scala 235:34]
  wire  _GEN_598 = ~io_inputBit | _GEN_597; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_599 = _GEN_6085 == 10'h241 ? _GEN_598 : _GEN_597; // @[lut_mem_online.scala 235:34]
  wire  _GEN_600 = io_inputBit ? 1'h0 : _GEN_599; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_601 = _GEN_6085 == 10'h241 ? _GEN_600 : _GEN_599; // @[lut_mem_online.scala 235:34]
  wire  _GEN_602 = ~io_inputBit ? 1'h0 : _GEN_601; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_603 = _GEN_6085 == 10'h242 ? _GEN_602 : _GEN_601; // @[lut_mem_online.scala 235:34]
  wire  _GEN_604 = io_inputBit | _GEN_603; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_605 = _GEN_6085 == 10'h242 ? _GEN_604 : _GEN_603; // @[lut_mem_online.scala 235:34]
  wire  _GEN_606 = ~io_inputBit | _GEN_605; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_607 = _GEN_6085 == 10'h243 ? _GEN_606 : _GEN_605; // @[lut_mem_online.scala 235:34]
  wire  _GEN_608 = io_inputBit ? 1'h0 : _GEN_607; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_609 = _GEN_6085 == 10'h243 ? _GEN_608 : _GEN_607; // @[lut_mem_online.scala 235:34]
  wire  _GEN_610 = ~io_inputBit ? 1'h0 : _GEN_609; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_611 = _GEN_6085 == 10'h244 ? _GEN_610 : _GEN_609; // @[lut_mem_online.scala 235:34]
  wire  _GEN_612 = io_inputBit | _GEN_611; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_613 = _GEN_6085 == 10'h244 ? _GEN_612 : _GEN_611; // @[lut_mem_online.scala 235:34]
  wire  _GEN_614 = ~io_inputBit | _GEN_613; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_615 = _GEN_6085 == 10'h245 ? _GEN_614 : _GEN_613; // @[lut_mem_online.scala 235:34]
  wire  _GEN_616 = io_inputBit ? 1'h0 : _GEN_615; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_617 = _GEN_6085 == 10'h245 ? _GEN_616 : _GEN_615; // @[lut_mem_online.scala 235:34]
  wire  _GEN_618 = ~io_inputBit ? 1'h0 : _GEN_617; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_619 = _GEN_6085 == 10'h246 ? _GEN_618 : _GEN_617; // @[lut_mem_online.scala 235:34]
  wire  _GEN_620 = io_inputBit | _GEN_619; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_621 = _GEN_6085 == 10'h246 ? _GEN_620 : _GEN_619; // @[lut_mem_online.scala 235:34]
  wire  _GEN_622 = ~io_inputBit | _GEN_621; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_623 = _GEN_6085 == 10'h247 ? _GEN_622 : _GEN_621; // @[lut_mem_online.scala 235:34]
  wire  _GEN_624 = io_inputBit ? 1'h0 : _GEN_623; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_625 = _GEN_6085 == 10'h247 ? _GEN_624 : _GEN_623; // @[lut_mem_online.scala 235:34]
  wire  _GEN_626 = ~io_inputBit ? 1'h0 : _GEN_625; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_627 = _GEN_6085 == 10'h248 ? _GEN_626 : _GEN_625; // @[lut_mem_online.scala 235:34]
  wire  _GEN_628 = io_inputBit | _GEN_627; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_629 = _GEN_6085 == 10'h248 ? _GEN_628 : _GEN_627; // @[lut_mem_online.scala 235:34]
  wire  _GEN_630 = ~io_inputBit | _GEN_629; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_631 = _GEN_6085 == 10'h249 ? _GEN_630 : _GEN_629; // @[lut_mem_online.scala 235:34]
  wire  _GEN_632 = io_inputBit ? 1'h0 : _GEN_631; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_633 = _GEN_6085 == 10'h249 ? _GEN_632 : _GEN_631; // @[lut_mem_online.scala 235:34]
  wire  _GEN_634 = io_inputBit ? 1'h0 : buffer_6; // @[lut_mem_online.scala 210:19 237:46 239:32]
  wire  _GEN_635 = i == 8'h0 ? _GEN_634 : buffer_6; // @[lut_mem_online.scala 210:19 235:34]
  wire  _GEN_636 = io_inputBit ? 1'h0 : _GEN_635; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_637 = i == 8'h1 ? _GEN_636 : _GEN_635; // @[lut_mem_online.scala 235:34]
  wire  _GEN_638 = io_inputBit ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_639 = i == 8'h8 ? _GEN_638 : _GEN_637; // @[lut_mem_online.scala 235:34]
  wire  _GEN_640 = ~io_inputBit ? 1'h0 : _GEN_639; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_641 = i == 8'hf ? _GEN_640 : _GEN_639; // @[lut_mem_online.scala 235:34]
  wire  _GEN_642 = io_inputBit ? 1'h0 : _GEN_641; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_643 = i == 8'h11 ? _GEN_642 : _GEN_641; // @[lut_mem_online.scala 235:34]
  wire  _GEN_644 = ~io_inputBit ? 1'h0 : _GEN_643; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_645 = i == 8'h20 ? _GEN_644 : _GEN_643; // @[lut_mem_online.scala 235:34]
  wire  _GEN_646 = io_inputBit ? 1'h0 : _GEN_645; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_647 = i == 8'h48 ? _GEN_646 : _GEN_645; // @[lut_mem_online.scala 235:34]
  wire  _GEN_648 = ~io_inputBit ? 1'h0 : _GEN_647; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_649 = _GEN_6084 == 9'h10b ? _GEN_648 : _GEN_647; // @[lut_mem_online.scala 235:34]
  wire  _GEN_650 = io_inputBit ? 1'h0 : _GEN_649; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_651 = _GEN_6084 == 9'h124 ? _GEN_650 : _GEN_649; // @[lut_mem_online.scala 235:34]
  wire  _GEN_652 = ~io_inputBit ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_653 = _GEN_6085 == 10'h218 ? _GEN_652 : _GEN_651; // @[lut_mem_online.scala 235:34]
  wire  _GEN_654 = io_inputBit | _GEN_653; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_655 = _GEN_6085 == 10'h218 ? _GEN_654 : _GEN_653; // @[lut_mem_online.scala 235:34]
  wire  _GEN_656 = ~io_inputBit ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_657 = _GEN_6085 == 10'h219 ? _GEN_656 : _GEN_655; // @[lut_mem_online.scala 235:34]
  wire  _GEN_658 = io_inputBit | _GEN_657; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_659 = _GEN_6085 == 10'h219 ? _GEN_658 : _GEN_657; // @[lut_mem_online.scala 235:34]
  wire  _GEN_660 = ~io_inputBit ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_661 = _GEN_6085 == 10'h21a ? _GEN_660 : _GEN_659; // @[lut_mem_online.scala 235:34]
  wire  _GEN_662 = io_inputBit | _GEN_661; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_663 = _GEN_6085 == 10'h21a ? _GEN_662 : _GEN_661; // @[lut_mem_online.scala 235:34]
  wire  _GEN_664 = ~io_inputBit ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_665 = _GEN_6085 == 10'h21b ? _GEN_664 : _GEN_663; // @[lut_mem_online.scala 235:34]
  wire  _GEN_666 = io_inputBit | _GEN_665; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_667 = _GEN_6085 == 10'h21b ? _GEN_666 : _GEN_665; // @[lut_mem_online.scala 235:34]
  wire  _GEN_668 = ~io_inputBit ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_669 = _GEN_6085 == 10'h21c ? _GEN_668 : _GEN_667; // @[lut_mem_online.scala 235:34]
  wire  _GEN_670 = io_inputBit | _GEN_669; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_671 = _GEN_6085 == 10'h21c ? _GEN_670 : _GEN_669; // @[lut_mem_online.scala 235:34]
  wire  _GEN_672 = ~io_inputBit ? 1'h0 : _GEN_671; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_673 = _GEN_6085 == 10'h21d ? _GEN_672 : _GEN_671; // @[lut_mem_online.scala 235:34]
  wire  _GEN_674 = io_inputBit | _GEN_673; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_675 = _GEN_6085 == 10'h21d ? _GEN_674 : _GEN_673; // @[lut_mem_online.scala 235:34]
  wire  _GEN_676 = ~io_inputBit ? 1'h0 : _GEN_675; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_677 = _GEN_6085 == 10'h21e ? _GEN_676 : _GEN_675; // @[lut_mem_online.scala 235:34]
  wire  _GEN_678 = io_inputBit | _GEN_677; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_679 = _GEN_6085 == 10'h21e ? _GEN_678 : _GEN_677; // @[lut_mem_online.scala 235:34]
  wire  _GEN_680 = ~io_inputBit ? 1'h0 : _GEN_679; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_681 = _GEN_6085 == 10'h21f ? _GEN_680 : _GEN_679; // @[lut_mem_online.scala 235:34]
  wire  _GEN_682 = io_inputBit | _GEN_681; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_683 = _GEN_6085 == 10'h21f ? _GEN_682 : _GEN_681; // @[lut_mem_online.scala 235:34]
  wire  _GEN_684 = ~io_inputBit ? 1'h0 : _GEN_683; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_685 = _GEN_6085 == 10'h220 ? _GEN_684 : _GEN_683; // @[lut_mem_online.scala 235:34]
  wire  _GEN_686 = io_inputBit | _GEN_685; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_687 = _GEN_6085 == 10'h220 ? _GEN_686 : _GEN_685; // @[lut_mem_online.scala 235:34]
  wire  _GEN_688 = ~io_inputBit ? 1'h0 : _GEN_687; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_689 = _GEN_6085 == 10'h221 ? _GEN_688 : _GEN_687; // @[lut_mem_online.scala 235:34]
  wire  _GEN_690 = io_inputBit | _GEN_689; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_691 = _GEN_6085 == 10'h221 ? _GEN_690 : _GEN_689; // @[lut_mem_online.scala 235:34]
  wire  _GEN_692 = ~io_inputBit ? 1'h0 : _GEN_691; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_693 = _GEN_6085 == 10'h222 ? _GEN_692 : _GEN_691; // @[lut_mem_online.scala 235:34]
  wire  _GEN_694 = io_inputBit | _GEN_693; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_695 = _GEN_6085 == 10'h222 ? _GEN_694 : _GEN_693; // @[lut_mem_online.scala 235:34]
  wire  _GEN_696 = ~io_inputBit ? 1'h0 : _GEN_695; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_697 = _GEN_6085 == 10'h223 ? _GEN_696 : _GEN_695; // @[lut_mem_online.scala 235:34]
  wire  _GEN_698 = io_inputBit | _GEN_697; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_699 = _GEN_6085 == 10'h223 ? _GEN_698 : _GEN_697; // @[lut_mem_online.scala 235:34]
  wire  _GEN_700 = ~io_inputBit ? 1'h0 : _GEN_699; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_701 = _GEN_6085 == 10'h224 ? _GEN_700 : _GEN_699; // @[lut_mem_online.scala 235:34]
  wire  _GEN_702 = io_inputBit | _GEN_701; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_703 = _GEN_6085 == 10'h224 ? _GEN_702 : _GEN_701; // @[lut_mem_online.scala 235:34]
  wire  _GEN_704 = ~io_inputBit ? 1'h0 : _GEN_703; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_705 = _GEN_6085 == 10'h225 ? _GEN_704 : _GEN_703; // @[lut_mem_online.scala 235:34]
  wire  _GEN_706 = io_inputBit | _GEN_705; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_707 = _GEN_6085 == 10'h225 ? _GEN_706 : _GEN_705; // @[lut_mem_online.scala 235:34]
  wire  _GEN_708 = ~io_inputBit ? 1'h0 : _GEN_707; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_709 = _GEN_6085 == 10'h226 ? _GEN_708 : _GEN_707; // @[lut_mem_online.scala 235:34]
  wire  _GEN_710 = io_inputBit | _GEN_709; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_711 = _GEN_6085 == 10'h226 ? _GEN_710 : _GEN_709; // @[lut_mem_online.scala 235:34]
  wire  _GEN_712 = ~io_inputBit ? 1'h0 : _GEN_711; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_713 = _GEN_6085 == 10'h227 ? _GEN_712 : _GEN_711; // @[lut_mem_online.scala 235:34]
  wire  _GEN_714 = io_inputBit | _GEN_713; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_715 = _GEN_6085 == 10'h227 ? _GEN_714 : _GEN_713; // @[lut_mem_online.scala 235:34]
  wire  _GEN_716 = ~io_inputBit ? 1'h0 : _GEN_715; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_717 = _GEN_6085 == 10'h228 ? _GEN_716 : _GEN_715; // @[lut_mem_online.scala 235:34]
  wire  _GEN_718 = io_inputBit | _GEN_717; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_719 = _GEN_6085 == 10'h228 ? _GEN_718 : _GEN_717; // @[lut_mem_online.scala 235:34]
  wire  _GEN_720 = ~io_inputBit ? 1'h0 : _GEN_719; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_721 = _GEN_6085 == 10'h229 ? _GEN_720 : _GEN_719; // @[lut_mem_online.scala 235:34]
  wire  _GEN_722 = io_inputBit | _GEN_721; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_723 = _GEN_6085 == 10'h229 ? _GEN_722 : _GEN_721; // @[lut_mem_online.scala 235:34]
  wire  _GEN_724 = ~io_inputBit ? 1'h0 : _GEN_723; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_725 = _GEN_6085 == 10'h22a ? _GEN_724 : _GEN_723; // @[lut_mem_online.scala 235:34]
  wire  _GEN_726 = io_inputBit | _GEN_725; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_727 = _GEN_6085 == 10'h22a ? _GEN_726 : _GEN_725; // @[lut_mem_online.scala 235:34]
  wire  _GEN_728 = ~io_inputBit ? 1'h0 : _GEN_727; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_729 = _GEN_6085 == 10'h22b ? _GEN_728 : _GEN_727; // @[lut_mem_online.scala 235:34]
  wire  _GEN_730 = io_inputBit | _GEN_729; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_731 = _GEN_6085 == 10'h22b ? _GEN_730 : _GEN_729; // @[lut_mem_online.scala 235:34]
  wire  _GEN_732 = ~io_inputBit ? 1'h0 : _GEN_731; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_733 = _GEN_6085 == 10'h22c ? _GEN_732 : _GEN_731; // @[lut_mem_online.scala 235:34]
  wire  _GEN_734 = io_inputBit | _GEN_733; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_735 = _GEN_6085 == 10'h22c ? _GEN_734 : _GEN_733; // @[lut_mem_online.scala 235:34]
  wire  _GEN_736 = ~io_inputBit ? 1'h0 : _GEN_735; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_737 = _GEN_6085 == 10'h22d ? _GEN_736 : _GEN_735; // @[lut_mem_online.scala 235:34]
  wire  _GEN_738 = io_inputBit | _GEN_737; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_739 = _GEN_6085 == 10'h22d ? _GEN_738 : _GEN_737; // @[lut_mem_online.scala 235:34]
  wire  _GEN_740 = ~io_inputBit ? 1'h0 : _GEN_739; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_741 = _GEN_6085 == 10'h22e ? _GEN_740 : _GEN_739; // @[lut_mem_online.scala 235:34]
  wire  _GEN_742 = io_inputBit | _GEN_741; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_743 = _GEN_6085 == 10'h22e ? _GEN_742 : _GEN_741; // @[lut_mem_online.scala 235:34]
  wire  _GEN_744 = ~io_inputBit ? 1'h0 : _GEN_743; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_745 = _GEN_6085 == 10'h22f ? _GEN_744 : _GEN_743; // @[lut_mem_online.scala 235:34]
  wire  _GEN_746 = io_inputBit | _GEN_745; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_747 = _GEN_6085 == 10'h22f ? _GEN_746 : _GEN_745; // @[lut_mem_online.scala 235:34]
  wire  _GEN_748 = ~io_inputBit ? 1'h0 : _GEN_747; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_749 = _GEN_6085 == 10'h230 ? _GEN_748 : _GEN_747; // @[lut_mem_online.scala 235:34]
  wire  _GEN_750 = io_inputBit | _GEN_749; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_751 = _GEN_6085 == 10'h230 ? _GEN_750 : _GEN_749; // @[lut_mem_online.scala 235:34]
  wire  _GEN_752 = ~io_inputBit ? 1'h0 : _GEN_751; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_753 = _GEN_6085 == 10'h231 ? _GEN_752 : _GEN_751; // @[lut_mem_online.scala 235:34]
  wire  _GEN_754 = io_inputBit | _GEN_753; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_755 = _GEN_6085 == 10'h231 ? _GEN_754 : _GEN_753; // @[lut_mem_online.scala 235:34]
  wire  _GEN_756 = ~io_inputBit ? 1'h0 : _GEN_755; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_757 = _GEN_6085 == 10'h232 ? _GEN_756 : _GEN_755; // @[lut_mem_online.scala 235:34]
  wire  _GEN_758 = io_inputBit | _GEN_757; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_759 = _GEN_6085 == 10'h232 ? _GEN_758 : _GEN_757; // @[lut_mem_online.scala 235:34]
  wire  _GEN_760 = ~io_inputBit ? 1'h0 : _GEN_759; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_761 = _GEN_6085 == 10'h233 ? _GEN_760 : _GEN_759; // @[lut_mem_online.scala 235:34]
  wire  _GEN_762 = io_inputBit | _GEN_761; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_763 = _GEN_6085 == 10'h233 ? _GEN_762 : _GEN_761; // @[lut_mem_online.scala 235:34]
  wire  _GEN_764 = ~io_inputBit ? 1'h0 : _GEN_763; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_765 = _GEN_6085 == 10'h234 ? _GEN_764 : _GEN_763; // @[lut_mem_online.scala 235:34]
  wire  _GEN_766 = io_inputBit | _GEN_765; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_767 = _GEN_6085 == 10'h234 ? _GEN_766 : _GEN_765; // @[lut_mem_online.scala 235:34]
  wire  _GEN_768 = ~io_inputBit ? 1'h0 : _GEN_767; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_769 = _GEN_6085 == 10'h235 ? _GEN_768 : _GEN_767; // @[lut_mem_online.scala 235:34]
  wire  _GEN_770 = io_inputBit | _GEN_769; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_771 = _GEN_6085 == 10'h235 ? _GEN_770 : _GEN_769; // @[lut_mem_online.scala 235:34]
  wire  _GEN_772 = ~io_inputBit ? 1'h0 : _GEN_771; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_773 = _GEN_6085 == 10'h236 ? _GEN_772 : _GEN_771; // @[lut_mem_online.scala 235:34]
  wire  _GEN_774 = io_inputBit | _GEN_773; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_775 = _GEN_6085 == 10'h236 ? _GEN_774 : _GEN_773; // @[lut_mem_online.scala 235:34]
  wire  _GEN_776 = ~io_inputBit ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_777 = _GEN_6085 == 10'h237 ? _GEN_776 : _GEN_775; // @[lut_mem_online.scala 235:34]
  wire  _GEN_778 = io_inputBit | _GEN_777; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_779 = _GEN_6085 == 10'h237 ? _GEN_778 : _GEN_777; // @[lut_mem_online.scala 235:34]
  wire  _GEN_780 = ~io_inputBit ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_781 = _GEN_6085 == 10'h238 ? _GEN_780 : _GEN_779; // @[lut_mem_online.scala 235:34]
  wire  _GEN_782 = io_inputBit | _GEN_781; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_783 = _GEN_6085 == 10'h238 ? _GEN_782 : _GEN_781; // @[lut_mem_online.scala 235:34]
  wire  _GEN_784 = ~io_inputBit ? 1'h0 : _GEN_783; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_785 = _GEN_6085 == 10'h239 ? _GEN_784 : _GEN_783; // @[lut_mem_online.scala 235:34]
  wire  _GEN_786 = io_inputBit | _GEN_785; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_787 = _GEN_6085 == 10'h239 ? _GEN_786 : _GEN_785; // @[lut_mem_online.scala 235:34]
  wire  _GEN_788 = ~io_inputBit ? 1'h0 : _GEN_787; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_789 = _GEN_6085 == 10'h23a ? _GEN_788 : _GEN_787; // @[lut_mem_online.scala 235:34]
  wire  _GEN_790 = io_inputBit | _GEN_789; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_791 = _GEN_6085 == 10'h23a ? _GEN_790 : _GEN_789; // @[lut_mem_online.scala 235:34]
  wire  _GEN_792 = ~io_inputBit ? 1'h0 : _GEN_791; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_793 = _GEN_6085 == 10'h23b ? _GEN_792 : _GEN_791; // @[lut_mem_online.scala 235:34]
  wire  _GEN_794 = io_inputBit | _GEN_793; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_795 = _GEN_6085 == 10'h23b ? _GEN_794 : _GEN_793; // @[lut_mem_online.scala 235:34]
  wire  _GEN_796 = ~io_inputBit ? 1'h0 : _GEN_795; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_797 = _GEN_6085 == 10'h23c ? _GEN_796 : _GEN_795; // @[lut_mem_online.scala 235:34]
  wire  _GEN_798 = io_inputBit | _GEN_797; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_799 = _GEN_6085 == 10'h23c ? _GEN_798 : _GEN_797; // @[lut_mem_online.scala 235:34]
  wire  _GEN_800 = ~io_inputBit ? 1'h0 : _GEN_799; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_801 = _GEN_6085 == 10'h23d ? _GEN_800 : _GEN_799; // @[lut_mem_online.scala 235:34]
  wire  _GEN_802 = io_inputBit | _GEN_801; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_803 = _GEN_6085 == 10'h23d ? _GEN_802 : _GEN_801; // @[lut_mem_online.scala 235:34]
  wire  _GEN_804 = ~io_inputBit ? 1'h0 : _GEN_803; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_805 = _GEN_6085 == 10'h23e ? _GEN_804 : _GEN_803; // @[lut_mem_online.scala 235:34]
  wire  _GEN_806 = io_inputBit | _GEN_805; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_807 = _GEN_6085 == 10'h23e ? _GEN_806 : _GEN_805; // @[lut_mem_online.scala 235:34]
  wire  _GEN_808 = ~io_inputBit ? 1'h0 : _GEN_807; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_809 = _GEN_6085 == 10'h23f ? _GEN_808 : _GEN_807; // @[lut_mem_online.scala 235:34]
  wire  _GEN_810 = io_inputBit | _GEN_809; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_811 = _GEN_6085 == 10'h23f ? _GEN_810 : _GEN_809; // @[lut_mem_online.scala 235:34]
  wire  _GEN_812 = ~io_inputBit ? 1'h0 : _GEN_811; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_813 = _GEN_6085 == 10'h240 ? _GEN_812 : _GEN_811; // @[lut_mem_online.scala 235:34]
  wire  _GEN_814 = io_inputBit | _GEN_813; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_815 = _GEN_6085 == 10'h240 ? _GEN_814 : _GEN_813; // @[lut_mem_online.scala 235:34]
  wire  _GEN_816 = ~io_inputBit ? 1'h0 : _GEN_815; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_817 = _GEN_6085 == 10'h241 ? _GEN_816 : _GEN_815; // @[lut_mem_online.scala 235:34]
  wire  _GEN_818 = io_inputBit | _GEN_817; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_819 = _GEN_6085 == 10'h241 ? _GEN_818 : _GEN_817; // @[lut_mem_online.scala 235:34]
  wire  _GEN_820 = ~io_inputBit ? 1'h0 : _GEN_819; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_821 = _GEN_6085 == 10'h242 ? _GEN_820 : _GEN_819; // @[lut_mem_online.scala 235:34]
  wire  _GEN_822 = io_inputBit | _GEN_821; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_823 = _GEN_6085 == 10'h242 ? _GEN_822 : _GEN_821; // @[lut_mem_online.scala 235:34]
  wire  _GEN_824 = ~io_inputBit ? 1'h0 : _GEN_823; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_825 = _GEN_6085 == 10'h243 ? _GEN_824 : _GEN_823; // @[lut_mem_online.scala 235:34]
  wire  _GEN_826 = io_inputBit | _GEN_825; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_827 = _GEN_6085 == 10'h243 ? _GEN_826 : _GEN_825; // @[lut_mem_online.scala 235:34]
  wire  _GEN_828 = ~io_inputBit ? 1'h0 : _GEN_827; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_829 = _GEN_6085 == 10'h244 ? _GEN_828 : _GEN_827; // @[lut_mem_online.scala 235:34]
  wire  _GEN_830 = io_inputBit | _GEN_829; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_831 = _GEN_6085 == 10'h244 ? _GEN_830 : _GEN_829; // @[lut_mem_online.scala 235:34]
  wire  _GEN_832 = ~io_inputBit ? 1'h0 : _GEN_831; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_833 = _GEN_6085 == 10'h245 ? _GEN_832 : _GEN_831; // @[lut_mem_online.scala 235:34]
  wire  _GEN_834 = io_inputBit | _GEN_833; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_835 = _GEN_6085 == 10'h245 ? _GEN_834 : _GEN_833; // @[lut_mem_online.scala 235:34]
  wire  _GEN_836 = ~io_inputBit ? 1'h0 : _GEN_835; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_837 = _GEN_6085 == 10'h246 ? _GEN_836 : _GEN_835; // @[lut_mem_online.scala 235:34]
  wire  _GEN_838 = io_inputBit | _GEN_837; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_839 = _GEN_6085 == 10'h246 ? _GEN_838 : _GEN_837; // @[lut_mem_online.scala 235:34]
  wire  _GEN_840 = ~io_inputBit ? 1'h0 : _GEN_839; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_841 = _GEN_6085 == 10'h247 ? _GEN_840 : _GEN_839; // @[lut_mem_online.scala 235:34]
  wire  _GEN_842 = io_inputBit | _GEN_841; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_843 = _GEN_6085 == 10'h247 ? _GEN_842 : _GEN_841; // @[lut_mem_online.scala 235:34]
  wire  _GEN_844 = ~io_inputBit ? 1'h0 : _GEN_843; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_845 = _GEN_6085 == 10'h248 ? _GEN_844 : _GEN_843; // @[lut_mem_online.scala 235:34]
  wire  _GEN_846 = io_inputBit | _GEN_845; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_847 = _GEN_6085 == 10'h248 ? _GEN_846 : _GEN_845; // @[lut_mem_online.scala 235:34]
  wire  _GEN_848 = ~io_inputBit ? 1'h0 : _GEN_847; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_849 = _GEN_6085 == 10'h249 ? _GEN_848 : _GEN_847; // @[lut_mem_online.scala 235:34]
  wire  _GEN_850 = io_inputBit | _GEN_849; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_851 = _GEN_6085 == 10'h249 ? _GEN_850 : _GEN_849; // @[lut_mem_online.scala 235:34]
  wire  _GEN_852 = io_inputBit ? 1'h0 : _GEN_21; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_853 = i == 8'h0 ? _GEN_852 : _GEN_21; // @[lut_mem_online.scala 235:34]
  wire  _GEN_854 = io_inputBit ? 1'h0 : _GEN_853; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_855 = i == 8'h1 ? _GEN_854 : _GEN_853; // @[lut_mem_online.scala 235:34]
  wire  _GEN_856 = ~io_inputBit ? 1'h0 : _GEN_855; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_857 = i == 8'h7 ? _GEN_856 : _GEN_855; // @[lut_mem_online.scala 235:34]
  wire  _GEN_858 = ~io_inputBit | _GEN_857; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_859 = i == 8'h8 ? _GEN_858 : _GEN_857; // @[lut_mem_online.scala 235:34]
  wire  _GEN_860 = ~io_inputBit ? 1'h0 : _GEN_859; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_861 = i == 8'h10 ? _GEN_860 : _GEN_859; // @[lut_mem_online.scala 235:34]
  wire  _GEN_862 = ~io_inputBit | _GEN_861; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_863 = i == 8'h12 ? _GEN_862 : _GEN_861; // @[lut_mem_online.scala 235:34]
  wire  _GEN_864 = ~io_inputBit ? 1'h0 : _GEN_863; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_865 = i == 8'h22 ? _GEN_864 : _GEN_863; // @[lut_mem_online.scala 235:34]
  wire  _GEN_866 = io_inputBit ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_867 = i == 8'h26 ? _GEN_866 : _GEN_865; // @[lut_mem_online.scala 235:34]
  wire  _GEN_868 = io_inputBit | _GEN_867; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_869 = i == 8'h46 ? _GEN_868 : _GEN_867; // @[lut_mem_online.scala 235:34]
  wire  _GEN_870 = ~io_inputBit | _GEN_869; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_871 = i == 8'h4d ? _GEN_870 : _GEN_869; // @[lut_mem_online.scala 235:34]
  wire  _GEN_872 = io_inputBit | _GEN_871; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_873 = i == 8'h8d ? _GEN_872 : _GEN_871; // @[lut_mem_online.scala 235:34]
  wire  _GEN_874 = ~io_inputBit | _GEN_873; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_875 = i == 8'h9c ? _GEN_874 : _GEN_873; // @[lut_mem_online.scala 235:34]
  wire  _GEN_876 = ~io_inputBit ? 1'h0 : _GEN_875; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_877 = _GEN_6084 == 9'h11b ? _GEN_876 : _GEN_875; // @[lut_mem_online.scala 235:34]
  wire  _GEN_878 = io_inputBit | _GEN_877; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_879 = _GEN_6084 == 9'h11b ? _GEN_878 : _GEN_877; // @[lut_mem_online.scala 235:34]
  wire  _GEN_880 = io_inputBit ? 1'h0 : _GEN_879; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_881 = _GEN_6084 == 9'h13a ? _GEN_880 : _GEN_879; // @[lut_mem_online.scala 235:34]
  wire  _GEN_882 = ~io_inputBit | _GEN_881; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_883 = _GEN_6085 == 10'h275 ? _GEN_882 : _GEN_881; // @[lut_mem_online.scala 235:34]
  wire  _GEN_884 = io_inputBit ? 1'h0 : _GEN_883; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_885 = _GEN_6085 == 10'h275 ? _GEN_884 : _GEN_883; // @[lut_mem_online.scala 235:34]
  wire  _GEN_886 = io_inputBit ? 1'h0 : _GEN_65; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_887 = i == 8'h0 ? _GEN_886 : _GEN_65; // @[lut_mem_online.scala 235:34]
  wire  _GEN_888 = io_inputBit ? 1'h0 : _GEN_887; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_889 = i == 8'h4 ? _GEN_888 : _GEN_887; // @[lut_mem_online.scala 235:34]
  wire  _GEN_890 = ~io_inputBit ? 1'h0 : _GEN_889; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_891 = i == 8'h7 ? _GEN_890 : _GEN_889; // @[lut_mem_online.scala 235:34]
  wire  _GEN_892 = io_inputBit ? 1'h0 : _GEN_891; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_893 = i == 8'h9 ? _GEN_892 : _GEN_891; // @[lut_mem_online.scala 235:34]
  wire  _GEN_894 = io_inputBit | _GEN_893; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_895 = i == 8'h11 ? _GEN_894 : _GEN_893; // @[lut_mem_online.scala 235:34]
  wire  _GEN_896 = io_inputBit ? 1'h0 : _GEN_895; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_897 = i == 8'h13 ? _GEN_896 : _GEN_895; // @[lut_mem_online.scala 235:34]
  wire  _GEN_898 = ~io_inputBit ? 1'h0 : _GEN_897; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_899 = i == 8'h21 ? _GEN_898 : _GEN_897; // @[lut_mem_online.scala 235:34]
  wire  _GEN_900 = ~io_inputBit | _GEN_899; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_901 = i == 8'h22 ? _GEN_900 : _GEN_899; // @[lut_mem_online.scala 235:34]
  wire  _GEN_902 = ~io_inputBit ? 1'h0 : _GEN_901; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_903 = i == 8'h23 ? _GEN_902 : _GEN_901; // @[lut_mem_online.scala 235:34]
  wire  _GEN_904 = io_inputBit ? 1'h0 : _GEN_903; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_905 = i == 8'h25 ? _GEN_904 : _GEN_903; // @[lut_mem_online.scala 235:34]
  wire  _GEN_906 = io_inputBit | _GEN_905; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_907 = i == 8'h26 ? _GEN_906 : _GEN_905; // @[lut_mem_online.scala 235:34]
  wire  _GEN_908 = io_inputBit ? 1'h0 : _GEN_907; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_909 = i == 8'h27 ? _GEN_908 : _GEN_907; // @[lut_mem_online.scala 235:34]
  wire  _GEN_910 = io_inputBit | _GEN_909; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_911 = i == 8'h44 ? _GEN_910 : _GEN_909; // @[lut_mem_online.scala 235:34]
  wire  _GEN_912 = io_inputBit ? 1'h0 : _GEN_911; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_913 = i == 8'h46 ? _GEN_912 : _GEN_911; // @[lut_mem_online.scala 235:34]
  wire  _GEN_914 = io_inputBit | _GEN_913; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_915 = i == 8'h48 ? _GEN_914 : _GEN_913; // @[lut_mem_online.scala 235:34]
  wire  _GEN_916 = ~io_inputBit | _GEN_915; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_917 = i == 8'h4b ? _GEN_916 : _GEN_915; // @[lut_mem_online.scala 235:34]
  wire  _GEN_918 = ~io_inputBit ? 1'h0 : _GEN_917; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_919 = i == 8'h4d ? _GEN_918 : _GEN_917; // @[lut_mem_online.scala 235:34]
  wire  _GEN_920 = ~io_inputBit | _GEN_919; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_921 = i == 8'h4f ? _GEN_920 : _GEN_919; // @[lut_mem_online.scala 235:34]
  wire  _GEN_922 = io_inputBit | _GEN_921; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_923 = i == 8'h89 ? _GEN_922 : _GEN_921; // @[lut_mem_online.scala 235:34]
  wire  _GEN_924 = io_inputBit ? 1'h0 : _GEN_923; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_925 = i == 8'h8d ? _GEN_924 : _GEN_923; // @[lut_mem_online.scala 235:34]
  wire  _GEN_926 = io_inputBit | _GEN_925; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_927 = i == 8'h91 ? _GEN_926 : _GEN_925; // @[lut_mem_online.scala 235:34]
  wire  _GEN_928 = ~io_inputBit | _GEN_927; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_929 = i == 8'h98 ? _GEN_928 : _GEN_927; // @[lut_mem_online.scala 235:34]
  wire  _GEN_930 = ~io_inputBit ? 1'h0 : _GEN_929; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_931 = i == 8'h9c ? _GEN_930 : _GEN_929; // @[lut_mem_online.scala 235:34]
  wire  _GEN_932 = ~io_inputBit | _GEN_931; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_933 = i == 8'ha0 ? _GEN_932 : _GEN_931; // @[lut_mem_online.scala 235:34]
  wire  _GEN_934 = ~io_inputBit ? 1'h0 : _GEN_933; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_935 = _GEN_6084 == 9'h113 ? _GEN_934 : _GEN_933; // @[lut_mem_online.scala 235:34]
  wire  _GEN_936 = io_inputBit | _GEN_935; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_937 = _GEN_6084 == 9'h113 ? _GEN_936 : _GEN_935; // @[lut_mem_online.scala 235:34]
  wire  _GEN_938 = ~io_inputBit | _GEN_937; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_939 = _GEN_6084 == 9'h11b ? _GEN_938 : _GEN_937; // @[lut_mem_online.scala 235:34]
  wire  _GEN_940 = io_inputBit ? 1'h0 : _GEN_939; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_941 = _GEN_6084 == 9'h11b ? _GEN_940 : _GEN_939; // @[lut_mem_online.scala 235:34]
  wire  _GEN_942 = ~io_inputBit ? 1'h0 : _GEN_941; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_943 = _GEN_6084 == 9'h123 ? _GEN_942 : _GEN_941; // @[lut_mem_online.scala 235:34]
  wire  _GEN_944 = io_inputBit | _GEN_943; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_945 = _GEN_6084 == 9'h123 ? _GEN_944 : _GEN_943; // @[lut_mem_online.scala 235:34]
  wire  _GEN_946 = io_inputBit ? 1'h0 : _GEN_945; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_947 = _GEN_6084 == 9'h132 ? _GEN_946 : _GEN_945; // @[lut_mem_online.scala 235:34]
  wire  _GEN_948 = io_inputBit | _GEN_947; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_949 = _GEN_6084 == 9'h13a ? _GEN_948 : _GEN_947; // @[lut_mem_online.scala 235:34]
  wire  _GEN_950 = io_inputBit ? 1'h0 : _GEN_949; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_951 = _GEN_6084 == 9'h142 ? _GEN_950 : _GEN_949; // @[lut_mem_online.scala 235:34]
  wire  _GEN_952 = ~io_inputBit | _GEN_951; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_953 = _GEN_6085 == 10'h265 ? _GEN_952 : _GEN_951; // @[lut_mem_online.scala 235:34]
  wire  _GEN_954 = io_inputBit ? 1'h0 : _GEN_953; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_955 = _GEN_6085 == 10'h265 ? _GEN_954 : _GEN_953; // @[lut_mem_online.scala 235:34]
  wire  _GEN_956 = ~io_inputBit ? 1'h0 : _GEN_955; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_957 = _GEN_6085 == 10'h275 ? _GEN_956 : _GEN_955; // @[lut_mem_online.scala 235:34]
  wire  _GEN_958 = io_inputBit | _GEN_957; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_959 = _GEN_6085 == 10'h275 ? _GEN_958 : _GEN_957; // @[lut_mem_online.scala 235:34]
  wire  _GEN_960 = ~io_inputBit | _GEN_959; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_961 = _GEN_6085 == 10'h285 ? _GEN_960 : _GEN_959; // @[lut_mem_online.scala 235:34]
  wire  _GEN_962 = io_inputBit ? 1'h0 : _GEN_961; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_963 = _GEN_6085 == 10'h285 ? _GEN_962 : _GEN_961; // @[lut_mem_online.scala 235:34]
  wire  _GEN_964 = io_inputBit ? 1'h0 : _GEN_139; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_965 = i == 8'h0 ? _GEN_964 : _GEN_139; // @[lut_mem_online.scala 235:34]
  wire  _GEN_966 = io_inputBit ? 1'h0 : _GEN_965; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_967 = i == 8'h4 ? _GEN_966 : _GEN_965; // @[lut_mem_online.scala 235:34]
  wire  _GEN_968 = ~io_inputBit ? 1'h0 : _GEN_967; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_969 = i == 8'h7 ? _GEN_968 : _GEN_967; // @[lut_mem_online.scala 235:34]
  wire  _GEN_970 = io_inputBit ? 1'h0 : _GEN_969; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_971 = i == 8'h9 ? _GEN_970 : _GEN_969; // @[lut_mem_online.scala 235:34]
  wire  _GEN_972 = io_inputBit ? 1'h0 : _GEN_971; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_973 = i == 8'h11 ? _GEN_972 : _GEN_971; // @[lut_mem_online.scala 235:34]
  wire  _GEN_974 = io_inputBit ? 1'h0 : _GEN_973; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_975 = i == 8'h13 ? _GEN_974 : _GEN_973; // @[lut_mem_online.scala 235:34]
  wire  _GEN_976 = io_inputBit | _GEN_975; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_977 = i == 8'h43 ? _GEN_976 : _GEN_975; // @[lut_mem_online.scala 235:34]
  wire  _GEN_978 = io_inputBit ? 1'h0 : _GEN_977; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_979 = i == 8'h44 ? _GEN_978 : _GEN_977; // @[lut_mem_online.scala 235:34]
  wire  _GEN_980 = io_inputBit | _GEN_979; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_981 = i == 8'h45 ? _GEN_980 : _GEN_979; // @[lut_mem_online.scala 235:34]
  wire  _GEN_982 = io_inputBit ? 1'h0 : _GEN_981; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_983 = i == 8'h46 ? _GEN_982 : _GEN_981; // @[lut_mem_online.scala 235:34]
  wire  _GEN_984 = io_inputBit | _GEN_983; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_985 = i == 8'h47 ? _GEN_984 : _GEN_983; // @[lut_mem_online.scala 235:34]
  wire  _GEN_986 = io_inputBit ? 1'h0 : _GEN_985; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_987 = i == 8'h48 ? _GEN_986 : _GEN_985; // @[lut_mem_online.scala 235:34]
  wire  _GEN_988 = ~io_inputBit ? 1'h0 : _GEN_987; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_989 = i == 8'h4b ? _GEN_988 : _GEN_987; // @[lut_mem_online.scala 235:34]
  wire  _GEN_990 = ~io_inputBit | _GEN_989; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_991 = i == 8'h4c ? _GEN_990 : _GEN_989; // @[lut_mem_online.scala 235:34]
  wire  _GEN_992 = ~io_inputBit ? 1'h0 : _GEN_991; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_993 = i == 8'h4d ? _GEN_992 : _GEN_991; // @[lut_mem_online.scala 235:34]
  wire  _GEN_994 = ~io_inputBit | _GEN_993; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_995 = i == 8'h4e ? _GEN_994 : _GEN_993; // @[lut_mem_online.scala 235:34]
  wire  _GEN_996 = ~io_inputBit ? 1'h0 : _GEN_995; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_997 = i == 8'h4f ? _GEN_996 : _GEN_995; // @[lut_mem_online.scala 235:34]
  wire  _GEN_998 = ~io_inputBit | _GEN_997; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_999 = i == 8'h50 ? _GEN_998 : _GEN_997; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1000 = io_inputBit | _GEN_999; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1001 = i == 8'h87 ? _GEN_1000 : _GEN_999; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1002 = io_inputBit ? 1'h0 : _GEN_1001; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1003 = i == 8'h89 ? _GEN_1002 : _GEN_1001; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1004 = io_inputBit | _GEN_1003; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1005 = i == 8'h8b ? _GEN_1004 : _GEN_1003; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1006 = io_inputBit ? 1'h0 : _GEN_1005; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1007 = i == 8'h8d ? _GEN_1006 : _GEN_1005; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1008 = io_inputBit | _GEN_1007; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1009 = i == 8'h8f ? _GEN_1008 : _GEN_1007; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1010 = io_inputBit ? 1'h0 : _GEN_1009; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1011 = i == 8'h91 ? _GEN_1010 : _GEN_1009; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1012 = ~io_inputBit ? 1'h0 : _GEN_1011; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1013 = i == 8'h98 ? _GEN_1012 : _GEN_1011; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1014 = ~io_inputBit | _GEN_1013; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1015 = i == 8'h9a ? _GEN_1014 : _GEN_1013; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1016 = ~io_inputBit ? 1'h0 : _GEN_1015; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1017 = i == 8'h9c ? _GEN_1016 : _GEN_1015; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1018 = ~io_inputBit | _GEN_1017; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1019 = i == 8'h9e ? _GEN_1018 : _GEN_1017; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1020 = ~io_inputBit ? 1'h0 : _GEN_1019; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1021 = i == 8'ha0 ? _GEN_1020 : _GEN_1019; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1022 = ~io_inputBit | _GEN_1021; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1023 = i == 8'ha2 ? _GEN_1022 : _GEN_1021; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1024 = ~io_inputBit ? 1'h0 : _GEN_1023; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1025 = _GEN_6084 == 9'h10f ? _GEN_1024 : _GEN_1023; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1026 = io_inputBit | _GEN_1025; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1027 = _GEN_6084 == 9'h10f ? _GEN_1026 : _GEN_1025; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1028 = ~io_inputBit | _GEN_1027; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1029 = _GEN_6084 == 9'h113 ? _GEN_1028 : _GEN_1027; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1030 = io_inputBit ? 1'h0 : _GEN_1029; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1031 = _GEN_6084 == 9'h113 ? _GEN_1030 : _GEN_1029; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1032 = ~io_inputBit ? 1'h0 : _GEN_1031; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1033 = _GEN_6084 == 9'h117 ? _GEN_1032 : _GEN_1031; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1034 = io_inputBit | _GEN_1033; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1035 = _GEN_6084 == 9'h117 ? _GEN_1034 : _GEN_1033; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1036 = ~io_inputBit | _GEN_1035; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1037 = _GEN_6084 == 9'h11b ? _GEN_1036 : _GEN_1035; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1038 = io_inputBit ? 1'h0 : _GEN_1037; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1039 = _GEN_6084 == 9'h11b ? _GEN_1038 : _GEN_1037; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1040 = ~io_inputBit ? 1'h0 : _GEN_1039; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1041 = _GEN_6084 == 9'h11f ? _GEN_1040 : _GEN_1039; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1042 = io_inputBit | _GEN_1041; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1043 = _GEN_6084 == 9'h11f ? _GEN_1042 : _GEN_1041; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1044 = ~io_inputBit | _GEN_1043; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1045 = _GEN_6084 == 9'h123 ? _GEN_1044 : _GEN_1043; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1046 = io_inputBit ? 1'h0 : _GEN_1045; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1047 = _GEN_6084 == 9'h123 ? _GEN_1046 : _GEN_1045; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1048 = io_inputBit | _GEN_1047; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1049 = _GEN_6084 == 9'h132 ? _GEN_1048 : _GEN_1047; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1050 = io_inputBit ? 1'h0 : _GEN_1049; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1051 = _GEN_6084 == 9'h136 ? _GEN_1050 : _GEN_1049; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1052 = io_inputBit | _GEN_1051; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1053 = _GEN_6084 == 9'h13a ? _GEN_1052 : _GEN_1051; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1054 = io_inputBit ? 1'h0 : _GEN_1053; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1055 = _GEN_6084 == 9'h13e ? _GEN_1054 : _GEN_1053; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1056 = io_inputBit | _GEN_1055; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1057 = _GEN_6084 == 9'h142 ? _GEN_1056 : _GEN_1055; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1058 = io_inputBit ? 1'h0 : _GEN_1057; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1059 = _GEN_6084 == 9'h146 ? _GEN_1058 : _GEN_1057; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1060 = ~io_inputBit ? 1'h0 : _GEN_1059; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1061 = _GEN_6085 == 10'h265 ? _GEN_1060 : _GEN_1059; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1062 = io_inputBit | _GEN_1061; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1063 = _GEN_6085 == 10'h265 ? _GEN_1062 : _GEN_1061; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1064 = ~io_inputBit | _GEN_1063; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1065 = _GEN_6085 == 10'h26d ? _GEN_1064 : _GEN_1063; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1066 = io_inputBit ? 1'h0 : _GEN_1065; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1067 = _GEN_6085 == 10'h26d ? _GEN_1066 : _GEN_1065; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1068 = ~io_inputBit ? 1'h0 : _GEN_1067; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1069 = _GEN_6085 == 10'h275 ? _GEN_1068 : _GEN_1067; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1070 = io_inputBit | _GEN_1069; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1071 = _GEN_6085 == 10'h275 ? _GEN_1070 : _GEN_1069; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1072 = ~io_inputBit | _GEN_1071; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1073 = _GEN_6085 == 10'h27d ? _GEN_1072 : _GEN_1071; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1074 = io_inputBit ? 1'h0 : _GEN_1073; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1075 = _GEN_6085 == 10'h27d ? _GEN_1074 : _GEN_1073; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1076 = ~io_inputBit ? 1'h0 : _GEN_1075; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1077 = _GEN_6085 == 10'h285 ? _GEN_1076 : _GEN_1075; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1078 = io_inputBit | _GEN_1077; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1079 = _GEN_6085 == 10'h285 ? _GEN_1078 : _GEN_1077; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1080 = ~io_inputBit | _GEN_1079; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1081 = _GEN_6085 == 10'h28d ? _GEN_1080 : _GEN_1079; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1082 = io_inputBit ? 1'h0 : _GEN_1081; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1083 = _GEN_6085 == 10'h28d ? _GEN_1082 : _GEN_1081; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1084 = io_inputBit ? 1'h0 : _GEN_249; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1085 = i == 8'h0 ? _GEN_1084 : _GEN_249; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1086 = io_inputBit ? 1'h0 : _GEN_1085; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1087 = i == 8'h4 ? _GEN_1086 : _GEN_1085; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1088 = io_inputBit ? 1'h0 : _GEN_1087; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1089 = i == 8'h9 ? _GEN_1088 : _GEN_1087; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1090 = ~io_inputBit ? 1'h0 : _GEN_1089; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1091 = i == 8'hf ? _GEN_1090 : _GEN_1089; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1092 = io_inputBit ? 1'h0 : _GEN_1091; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1093 = i == 8'h11 ? _GEN_1092 : _GEN_1091; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1094 = ~io_inputBit ? 1'h0 : _GEN_1093; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1095 = i == 8'h20 ? _GEN_1094 : _GEN_1093; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1096 = io_inputBit ? 1'h0 : _GEN_1095; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1097 = i == 8'h28 ? _GEN_1096 : _GEN_1095; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1098 = ~io_inputBit ? 1'h0 : _GEN_1097; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1099 = i == 8'h42 ? _GEN_1098 : _GEN_1097; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1100 = io_inputBit ? 1'h0 : _GEN_1099; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1101 = i == 8'h48 ? _GEN_1100 : _GEN_1099; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1102 = ~io_inputBit ? 1'h0 : _GEN_1101; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1103 = i == 8'h4b ? _GEN_1102 : _GEN_1101; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1104 = io_inputBit ? 1'h0 : _GEN_1103; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1105 = i == 8'h51 ? _GEN_1104 : _GEN_1103; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1106 = io_inputBit | _GEN_1105; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1107 = i == 8'h86 ? _GEN_1106 : _GEN_1105; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1108 = io_inputBit ? 1'h0 : _GEN_1107; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1109 = i == 8'h87 ? _GEN_1108 : _GEN_1107; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1110 = io_inputBit | _GEN_1109; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1111 = i == 8'h88 ? _GEN_1110 : _GEN_1109; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1112 = io_inputBit ? 1'h0 : _GEN_1111; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1113 = i == 8'h89 ? _GEN_1112 : _GEN_1111; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1114 = io_inputBit | _GEN_1113; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1115 = i == 8'h8a ? _GEN_1114 : _GEN_1113; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1116 = io_inputBit ? 1'h0 : _GEN_1115; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1117 = i == 8'h8b ? _GEN_1116 : _GEN_1115; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1118 = io_inputBit | _GEN_1117; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1119 = i == 8'h8c ? _GEN_1118 : _GEN_1117; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1120 = io_inputBit ? 1'h0 : _GEN_1119; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1121 = i == 8'h8d ? _GEN_1120 : _GEN_1119; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1122 = io_inputBit | _GEN_1121; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1123 = i == 8'h8e ? _GEN_1122 : _GEN_1121; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1124 = io_inputBit ? 1'h0 : _GEN_1123; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1125 = i == 8'h8f ? _GEN_1124 : _GEN_1123; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1126 = io_inputBit | _GEN_1125; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1127 = i == 8'h90 ? _GEN_1126 : _GEN_1125; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1128 = io_inputBit ? 1'h0 : _GEN_1127; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1129 = i == 8'h91 ? _GEN_1128 : _GEN_1127; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1130 = ~io_inputBit ? 1'h0 : _GEN_1129; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1131 = i == 8'h98 ? _GEN_1130 : _GEN_1129; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1132 = ~io_inputBit | _GEN_1131; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1133 = i == 8'h99 ? _GEN_1132 : _GEN_1131; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1134 = ~io_inputBit ? 1'h0 : _GEN_1133; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1135 = i == 8'h9a ? _GEN_1134 : _GEN_1133; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1136 = ~io_inputBit | _GEN_1135; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1137 = i == 8'h9b ? _GEN_1136 : _GEN_1135; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1138 = ~io_inputBit ? 1'h0 : _GEN_1137; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1139 = i == 8'h9c ? _GEN_1138 : _GEN_1137; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1140 = ~io_inputBit | _GEN_1139; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1141 = i == 8'h9d ? _GEN_1140 : _GEN_1139; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1142 = ~io_inputBit ? 1'h0 : _GEN_1141; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1143 = i == 8'h9e ? _GEN_1142 : _GEN_1141; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1144 = ~io_inputBit | _GEN_1143; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1145 = i == 8'h9f ? _GEN_1144 : _GEN_1143; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1146 = ~io_inputBit ? 1'h0 : _GEN_1145; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1147 = i == 8'ha0 ? _GEN_1146 : _GEN_1145; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1148 = ~io_inputBit | _GEN_1147; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1149 = i == 8'ha1 ? _GEN_1148 : _GEN_1147; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1150 = ~io_inputBit ? 1'h0 : _GEN_1149; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1151 = i == 8'ha2 ? _GEN_1150 : _GEN_1149; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1152 = ~io_inputBit | _GEN_1151; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1153 = i == 8'ha3 ? _GEN_1152 : _GEN_1151; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1154 = ~io_inputBit ? 1'h0 : _GEN_1153; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1155 = _GEN_6084 == 9'h10d ? _GEN_1154 : _GEN_1153; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1156 = io_inputBit | _GEN_1155; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1157 = _GEN_6084 == 9'h10d ? _GEN_1156 : _GEN_1155; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1158 = ~io_inputBit | _GEN_1157; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1159 = _GEN_6084 == 9'h10f ? _GEN_1158 : _GEN_1157; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1160 = io_inputBit ? 1'h0 : _GEN_1159; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1161 = _GEN_6084 == 9'h10f ? _GEN_1160 : _GEN_1159; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1162 = ~io_inputBit ? 1'h0 : _GEN_1161; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1163 = _GEN_6084 == 9'h111 ? _GEN_1162 : _GEN_1161; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1164 = io_inputBit | _GEN_1163; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1165 = _GEN_6084 == 9'h111 ? _GEN_1164 : _GEN_1163; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1166 = ~io_inputBit | _GEN_1165; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1167 = _GEN_6084 == 9'h113 ? _GEN_1166 : _GEN_1165; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1168 = io_inputBit ? 1'h0 : _GEN_1167; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1169 = _GEN_6084 == 9'h113 ? _GEN_1168 : _GEN_1167; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1170 = ~io_inputBit ? 1'h0 : _GEN_1169; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1171 = _GEN_6084 == 9'h115 ? _GEN_1170 : _GEN_1169; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1172 = io_inputBit | _GEN_1171; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1173 = _GEN_6084 == 9'h115 ? _GEN_1172 : _GEN_1171; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1174 = ~io_inputBit | _GEN_1173; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1175 = _GEN_6084 == 9'h117 ? _GEN_1174 : _GEN_1173; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1176 = io_inputBit ? 1'h0 : _GEN_1175; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1177 = _GEN_6084 == 9'h117 ? _GEN_1176 : _GEN_1175; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1178 = ~io_inputBit ? 1'h0 : _GEN_1177; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1179 = _GEN_6084 == 9'h119 ? _GEN_1178 : _GEN_1177; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1180 = io_inputBit | _GEN_1179; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1181 = _GEN_6084 == 9'h119 ? _GEN_1180 : _GEN_1179; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1182 = ~io_inputBit | _GEN_1181; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1183 = _GEN_6084 == 9'h11b ? _GEN_1182 : _GEN_1181; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1184 = io_inputBit ? 1'h0 : _GEN_1183; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1185 = _GEN_6084 == 9'h11b ? _GEN_1184 : _GEN_1183; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1186 = ~io_inputBit ? 1'h0 : _GEN_1185; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1187 = _GEN_6084 == 9'h11d ? _GEN_1186 : _GEN_1185; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1188 = io_inputBit | _GEN_1187; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1189 = _GEN_6084 == 9'h11d ? _GEN_1188 : _GEN_1187; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1190 = ~io_inputBit | _GEN_1189; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1191 = _GEN_6084 == 9'h11f ? _GEN_1190 : _GEN_1189; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1192 = io_inputBit ? 1'h0 : _GEN_1191; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1193 = _GEN_6084 == 9'h11f ? _GEN_1192 : _GEN_1191; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1194 = ~io_inputBit ? 1'h0 : _GEN_1193; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1195 = _GEN_6084 == 9'h121 ? _GEN_1194 : _GEN_1193; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1196 = io_inputBit | _GEN_1195; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1197 = _GEN_6084 == 9'h121 ? _GEN_1196 : _GEN_1195; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1198 = ~io_inputBit | _GEN_1197; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1199 = _GEN_6084 == 9'h123 ? _GEN_1198 : _GEN_1197; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1200 = io_inputBit ? 1'h0 : _GEN_1199; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1201 = _GEN_6084 == 9'h123 ? _GEN_1200 : _GEN_1199; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1202 = io_inputBit | _GEN_1201; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1203 = _GEN_6084 == 9'h132 ? _GEN_1202 : _GEN_1201; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1204 = io_inputBit ? 1'h0 : _GEN_1203; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1205 = _GEN_6084 == 9'h134 ? _GEN_1204 : _GEN_1203; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1206 = io_inputBit | _GEN_1205; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1207 = _GEN_6084 == 9'h136 ? _GEN_1206 : _GEN_1205; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1208 = io_inputBit ? 1'h0 : _GEN_1207; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1209 = _GEN_6084 == 9'h138 ? _GEN_1208 : _GEN_1207; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1210 = io_inputBit | _GEN_1209; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1211 = _GEN_6084 == 9'h13a ? _GEN_1210 : _GEN_1209; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1212 = io_inputBit ? 1'h0 : _GEN_1211; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1213 = _GEN_6084 == 9'h13c ? _GEN_1212 : _GEN_1211; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1214 = io_inputBit | _GEN_1213; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1215 = _GEN_6084 == 9'h13e ? _GEN_1214 : _GEN_1213; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1216 = io_inputBit ? 1'h0 : _GEN_1215; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1217 = _GEN_6084 == 9'h140 ? _GEN_1216 : _GEN_1215; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1218 = io_inputBit | _GEN_1217; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1219 = _GEN_6084 == 9'h142 ? _GEN_1218 : _GEN_1217; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1220 = io_inputBit ? 1'h0 : _GEN_1219; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1221 = _GEN_6084 == 9'h144 ? _GEN_1220 : _GEN_1219; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1222 = io_inputBit | _GEN_1221; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1223 = _GEN_6084 == 9'h146 ? _GEN_1222 : _GEN_1221; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1224 = io_inputBit ? 1'h0 : _GEN_1223; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1225 = _GEN_6084 == 9'h148 ? _GEN_1224 : _GEN_1223; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1226 = ~io_inputBit ? 1'h0 : _GEN_1225; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1227 = _GEN_6085 == 10'h265 ? _GEN_1226 : _GEN_1225; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1228 = io_inputBit | _GEN_1227; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1229 = _GEN_6085 == 10'h265 ? _GEN_1228 : _GEN_1227; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1230 = ~io_inputBit | _GEN_1229; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1231 = _GEN_6085 == 10'h269 ? _GEN_1230 : _GEN_1229; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1232 = io_inputBit ? 1'h0 : _GEN_1231; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1233 = _GEN_6085 == 10'h269 ? _GEN_1232 : _GEN_1231; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1234 = ~io_inputBit ? 1'h0 : _GEN_1233; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1235 = _GEN_6085 == 10'h26d ? _GEN_1234 : _GEN_1233; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1236 = io_inputBit | _GEN_1235; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1237 = _GEN_6085 == 10'h26d ? _GEN_1236 : _GEN_1235; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1238 = ~io_inputBit | _GEN_1237; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1239 = _GEN_6085 == 10'h271 ? _GEN_1238 : _GEN_1237; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1240 = io_inputBit ? 1'h0 : _GEN_1239; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1241 = _GEN_6085 == 10'h271 ? _GEN_1240 : _GEN_1239; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1242 = ~io_inputBit ? 1'h0 : _GEN_1241; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1243 = _GEN_6085 == 10'h275 ? _GEN_1242 : _GEN_1241; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1244 = io_inputBit | _GEN_1243; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1245 = _GEN_6085 == 10'h275 ? _GEN_1244 : _GEN_1243; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1246 = ~io_inputBit | _GEN_1245; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1247 = _GEN_6085 == 10'h279 ? _GEN_1246 : _GEN_1245; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1248 = io_inputBit ? 1'h0 : _GEN_1247; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1249 = _GEN_6085 == 10'h279 ? _GEN_1248 : _GEN_1247; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1250 = ~io_inputBit ? 1'h0 : _GEN_1249; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1251 = _GEN_6085 == 10'h27d ? _GEN_1250 : _GEN_1249; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1252 = io_inputBit | _GEN_1251; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1253 = _GEN_6085 == 10'h27d ? _GEN_1252 : _GEN_1251; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1254 = ~io_inputBit | _GEN_1253; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1255 = _GEN_6085 == 10'h281 ? _GEN_1254 : _GEN_1253; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1256 = io_inputBit ? 1'h0 : _GEN_1255; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1257 = _GEN_6085 == 10'h281 ? _GEN_1256 : _GEN_1255; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1258 = ~io_inputBit ? 1'h0 : _GEN_1257; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1259 = _GEN_6085 == 10'h285 ? _GEN_1258 : _GEN_1257; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1260 = io_inputBit | _GEN_1259; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1261 = _GEN_6085 == 10'h285 ? _GEN_1260 : _GEN_1259; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1262 = ~io_inputBit | _GEN_1261; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1263 = _GEN_6085 == 10'h289 ? _GEN_1262 : _GEN_1261; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1264 = io_inputBit ? 1'h0 : _GEN_1263; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1265 = _GEN_6085 == 10'h289 ? _GEN_1264 : _GEN_1263; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1266 = ~io_inputBit ? 1'h0 : _GEN_1265; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1267 = _GEN_6085 == 10'h28d ? _GEN_1266 : _GEN_1265; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1268 = io_inputBit | _GEN_1267; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1269 = _GEN_6085 == 10'h28d ? _GEN_1268 : _GEN_1267; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1270 = ~io_inputBit | _GEN_1269; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1271 = _GEN_6085 == 10'h291 ? _GEN_1270 : _GEN_1269; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1272 = io_inputBit ? 1'h0 : _GEN_1271; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1273 = _GEN_6085 == 10'h291 ? _GEN_1272 : _GEN_1271; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1274 = io_inputBit ? 1'h0 : _GEN_415; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1275 = i == 8'h0 ? _GEN_1274 : _GEN_415; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1276 = io_inputBit ? 1'h0 : _GEN_1275; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1277 = i == 8'h4 ? _GEN_1276 : _GEN_1275; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1278 = io_inputBit ? 1'h0 : _GEN_1277; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1279 = i == 8'h9 ? _GEN_1278 : _GEN_1277; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1280 = ~io_inputBit ? 1'h0 : _GEN_1279; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1281 = i == 8'hf ? _GEN_1280 : _GEN_1279; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1282 = io_inputBit | _GEN_1281; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1283 = i == 8'h11 ? _GEN_1282 : _GEN_1281; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1284 = ~io_inputBit ? 1'h0 : _GEN_1283; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1285 = i == 8'h20 ? _GEN_1284 : _GEN_1283; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1286 = io_inputBit ? 1'h0 : _GEN_1285; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1287 = i == 8'h28 ? _GEN_1286 : _GEN_1285; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1288 = io_inputBit | _GEN_1287; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1289 = i == 8'h48 ? _GEN_1288 : _GEN_1287; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1290 = ~io_inputBit | _GEN_1289; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1291 = i == 8'h4b ? _GEN_1290 : _GEN_1289; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1292 = ~io_inputBit ? 1'h0 : _GEN_1291; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1293 = i == 8'h85 ? _GEN_1292 : _GEN_1291; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1294 = io_inputBit ? 1'h0 : _GEN_1293; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1295 = i == 8'ha4 ? _GEN_1294 : _GEN_1293; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1296 = ~io_inputBit ? 1'h0 : _GEN_1295; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1297 = _GEN_6084 == 9'h10c ? _GEN_1296 : _GEN_1295; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1298 = io_inputBit | _GEN_1297; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1299 = _GEN_6084 == 9'h10c ? _GEN_1298 : _GEN_1297; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1300 = ~io_inputBit | _GEN_1299; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1301 = _GEN_6084 == 9'h10d ? _GEN_1300 : _GEN_1299; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1302 = io_inputBit ? 1'h0 : _GEN_1301; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1303 = _GEN_6084 == 9'h10d ? _GEN_1302 : _GEN_1301; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1304 = ~io_inputBit ? 1'h0 : _GEN_1303; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1305 = _GEN_6084 == 9'h10e ? _GEN_1304 : _GEN_1303; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1306 = io_inputBit | _GEN_1305; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1307 = _GEN_6084 == 9'h10e ? _GEN_1306 : _GEN_1305; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1308 = ~io_inputBit | _GEN_1307; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1309 = _GEN_6084 == 9'h10f ? _GEN_1308 : _GEN_1307; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1310 = io_inputBit ? 1'h0 : _GEN_1309; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1311 = _GEN_6084 == 9'h10f ? _GEN_1310 : _GEN_1309; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1312 = ~io_inputBit ? 1'h0 : _GEN_1311; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1313 = _GEN_6084 == 9'h110 ? _GEN_1312 : _GEN_1311; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1314 = io_inputBit | _GEN_1313; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1315 = _GEN_6084 == 9'h110 ? _GEN_1314 : _GEN_1313; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1316 = ~io_inputBit | _GEN_1315; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1317 = _GEN_6084 == 9'h111 ? _GEN_1316 : _GEN_1315; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1318 = io_inputBit ? 1'h0 : _GEN_1317; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1319 = _GEN_6084 == 9'h111 ? _GEN_1318 : _GEN_1317; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1320 = ~io_inputBit ? 1'h0 : _GEN_1319; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1321 = _GEN_6084 == 9'h112 ? _GEN_1320 : _GEN_1319; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1322 = io_inputBit | _GEN_1321; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1323 = _GEN_6084 == 9'h112 ? _GEN_1322 : _GEN_1321; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1324 = ~io_inputBit | _GEN_1323; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1325 = _GEN_6084 == 9'h113 ? _GEN_1324 : _GEN_1323; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1326 = io_inputBit ? 1'h0 : _GEN_1325; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1327 = _GEN_6084 == 9'h113 ? _GEN_1326 : _GEN_1325; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1328 = ~io_inputBit ? 1'h0 : _GEN_1327; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1329 = _GEN_6084 == 9'h114 ? _GEN_1328 : _GEN_1327; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1330 = io_inputBit | _GEN_1329; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1331 = _GEN_6084 == 9'h114 ? _GEN_1330 : _GEN_1329; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1332 = ~io_inputBit | _GEN_1331; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1333 = _GEN_6084 == 9'h115 ? _GEN_1332 : _GEN_1331; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1334 = io_inputBit ? 1'h0 : _GEN_1333; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1335 = _GEN_6084 == 9'h115 ? _GEN_1334 : _GEN_1333; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1336 = ~io_inputBit ? 1'h0 : _GEN_1335; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1337 = _GEN_6084 == 9'h116 ? _GEN_1336 : _GEN_1335; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1338 = io_inputBit | _GEN_1337; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1339 = _GEN_6084 == 9'h116 ? _GEN_1338 : _GEN_1337; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1340 = ~io_inputBit | _GEN_1339; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1341 = _GEN_6084 == 9'h117 ? _GEN_1340 : _GEN_1339; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1342 = io_inputBit ? 1'h0 : _GEN_1341; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1343 = _GEN_6084 == 9'h117 ? _GEN_1342 : _GEN_1341; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1344 = ~io_inputBit ? 1'h0 : _GEN_1343; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1345 = _GEN_6084 == 9'h118 ? _GEN_1344 : _GEN_1343; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1346 = io_inputBit | _GEN_1345; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1347 = _GEN_6084 == 9'h118 ? _GEN_1346 : _GEN_1345; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1348 = ~io_inputBit | _GEN_1347; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1349 = _GEN_6084 == 9'h119 ? _GEN_1348 : _GEN_1347; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1350 = io_inputBit ? 1'h0 : _GEN_1349; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1351 = _GEN_6084 == 9'h119 ? _GEN_1350 : _GEN_1349; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1352 = ~io_inputBit ? 1'h0 : _GEN_1351; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1353 = _GEN_6084 == 9'h11a ? _GEN_1352 : _GEN_1351; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1354 = io_inputBit | _GEN_1353; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1355 = _GEN_6084 == 9'h11a ? _GEN_1354 : _GEN_1353; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1356 = ~io_inputBit | _GEN_1355; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1357 = _GEN_6084 == 9'h11b ? _GEN_1356 : _GEN_1355; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1358 = io_inputBit ? 1'h0 : _GEN_1357; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1359 = _GEN_6084 == 9'h11b ? _GEN_1358 : _GEN_1357; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1360 = ~io_inputBit ? 1'h0 : _GEN_1359; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1361 = _GEN_6084 == 9'h11c ? _GEN_1360 : _GEN_1359; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1362 = io_inputBit | _GEN_1361; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1363 = _GEN_6084 == 9'h11c ? _GEN_1362 : _GEN_1361; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1364 = ~io_inputBit | _GEN_1363; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1365 = _GEN_6084 == 9'h11d ? _GEN_1364 : _GEN_1363; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1366 = io_inputBit ? 1'h0 : _GEN_1365; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1367 = _GEN_6084 == 9'h11d ? _GEN_1366 : _GEN_1365; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1368 = ~io_inputBit ? 1'h0 : _GEN_1367; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1369 = _GEN_6084 == 9'h11e ? _GEN_1368 : _GEN_1367; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1370 = io_inputBit | _GEN_1369; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1371 = _GEN_6084 == 9'h11e ? _GEN_1370 : _GEN_1369; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1372 = ~io_inputBit | _GEN_1371; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1373 = _GEN_6084 == 9'h11f ? _GEN_1372 : _GEN_1371; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1374 = io_inputBit ? 1'h0 : _GEN_1373; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1375 = _GEN_6084 == 9'h11f ? _GEN_1374 : _GEN_1373; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1376 = ~io_inputBit ? 1'h0 : _GEN_1375; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1377 = _GEN_6084 == 9'h120 ? _GEN_1376 : _GEN_1375; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1378 = io_inputBit | _GEN_1377; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1379 = _GEN_6084 == 9'h120 ? _GEN_1378 : _GEN_1377; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1380 = ~io_inputBit | _GEN_1379; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1381 = _GEN_6084 == 9'h121 ? _GEN_1380 : _GEN_1379; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1382 = io_inputBit ? 1'h0 : _GEN_1381; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1383 = _GEN_6084 == 9'h121 ? _GEN_1382 : _GEN_1381; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1384 = ~io_inputBit ? 1'h0 : _GEN_1383; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1385 = _GEN_6084 == 9'h122 ? _GEN_1384 : _GEN_1383; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1386 = io_inputBit | _GEN_1385; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1387 = _GEN_6084 == 9'h122 ? _GEN_1386 : _GEN_1385; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1388 = ~io_inputBit | _GEN_1387; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1389 = _GEN_6084 == 9'h123 ? _GEN_1388 : _GEN_1387; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1390 = io_inputBit ? 1'h0 : _GEN_1389; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1391 = _GEN_6084 == 9'h123 ? _GEN_1390 : _GEN_1389; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1392 = ~io_inputBit ? 1'h0 : _GEN_1391; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1393 = _GEN_6084 == 9'h124 ? _GEN_1392 : _GEN_1391; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1394 = io_inputBit | _GEN_1393; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1395 = _GEN_6084 == 9'h124 ? _GEN_1394 : _GEN_1393; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1396 = io_inputBit ? 1'h0 : _GEN_1395; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1397 = _GEN_6084 == 9'h131 ? _GEN_1396 : _GEN_1395; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1398 = io_inputBit | _GEN_1397; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1399 = _GEN_6084 == 9'h132 ? _GEN_1398 : _GEN_1397; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1400 = io_inputBit ? 1'h0 : _GEN_1399; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1401 = _GEN_6084 == 9'h133 ? _GEN_1400 : _GEN_1399; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1402 = io_inputBit | _GEN_1401; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1403 = _GEN_6084 == 9'h134 ? _GEN_1402 : _GEN_1401; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1404 = io_inputBit ? 1'h0 : _GEN_1403; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1405 = _GEN_6084 == 9'h135 ? _GEN_1404 : _GEN_1403; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1406 = io_inputBit | _GEN_1405; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1407 = _GEN_6084 == 9'h136 ? _GEN_1406 : _GEN_1405; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1408 = io_inputBit ? 1'h0 : _GEN_1407; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1409 = _GEN_6084 == 9'h137 ? _GEN_1408 : _GEN_1407; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1410 = io_inputBit | _GEN_1409; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1411 = _GEN_6084 == 9'h138 ? _GEN_1410 : _GEN_1409; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1412 = io_inputBit ? 1'h0 : _GEN_1411; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1413 = _GEN_6084 == 9'h139 ? _GEN_1412 : _GEN_1411; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1414 = io_inputBit | _GEN_1413; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1415 = _GEN_6084 == 9'h13a ? _GEN_1414 : _GEN_1413; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1416 = io_inputBit ? 1'h0 : _GEN_1415; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1417 = _GEN_6084 == 9'h13b ? _GEN_1416 : _GEN_1415; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1418 = io_inputBit | _GEN_1417; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1419 = _GEN_6084 == 9'h13c ? _GEN_1418 : _GEN_1417; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1420 = io_inputBit ? 1'h0 : _GEN_1419; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1421 = _GEN_6084 == 9'h13d ? _GEN_1420 : _GEN_1419; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1422 = io_inputBit | _GEN_1421; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1423 = _GEN_6084 == 9'h13e ? _GEN_1422 : _GEN_1421; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1424 = io_inputBit ? 1'h0 : _GEN_1423; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1425 = _GEN_6084 == 9'h13f ? _GEN_1424 : _GEN_1423; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1426 = io_inputBit | _GEN_1425; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1427 = _GEN_6084 == 9'h140 ? _GEN_1426 : _GEN_1425; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1428 = io_inputBit ? 1'h0 : _GEN_1427; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1429 = _GEN_6084 == 9'h141 ? _GEN_1428 : _GEN_1427; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1430 = io_inputBit | _GEN_1429; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1431 = _GEN_6084 == 9'h142 ? _GEN_1430 : _GEN_1429; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1432 = io_inputBit ? 1'h0 : _GEN_1431; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1433 = _GEN_6084 == 9'h143 ? _GEN_1432 : _GEN_1431; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1434 = io_inputBit | _GEN_1433; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1435 = _GEN_6084 == 9'h144 ? _GEN_1434 : _GEN_1433; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1436 = io_inputBit ? 1'h0 : _GEN_1435; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1437 = _GEN_6084 == 9'h145 ? _GEN_1436 : _GEN_1435; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1438 = io_inputBit | _GEN_1437; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1439 = _GEN_6084 == 9'h146 ? _GEN_1438 : _GEN_1437; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1440 = io_inputBit ? 1'h0 : _GEN_1439; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1441 = _GEN_6084 == 9'h147 ? _GEN_1440 : _GEN_1439; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1442 = io_inputBit | _GEN_1441; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1443 = _GEN_6084 == 9'h148 ? _GEN_1442 : _GEN_1441; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1444 = io_inputBit ? 1'h0 : _GEN_1443; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1445 = _GEN_6084 == 9'h149 ? _GEN_1444 : _GEN_1443; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1446 = ~io_inputBit | _GEN_1445; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1447 = _GEN_6085 == 10'h263 ? _GEN_1446 : _GEN_1445; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1448 = io_inputBit ? 1'h0 : _GEN_1447; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1449 = _GEN_6085 == 10'h263 ? _GEN_1448 : _GEN_1447; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1450 = ~io_inputBit ? 1'h0 : _GEN_1449; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1451 = _GEN_6085 == 10'h265 ? _GEN_1450 : _GEN_1449; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1452 = io_inputBit | _GEN_1451; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1453 = _GEN_6085 == 10'h265 ? _GEN_1452 : _GEN_1451; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1454 = ~io_inputBit | _GEN_1453; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1455 = _GEN_6085 == 10'h267 ? _GEN_1454 : _GEN_1453; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1456 = io_inputBit ? 1'h0 : _GEN_1455; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1457 = _GEN_6085 == 10'h267 ? _GEN_1456 : _GEN_1455; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1458 = ~io_inputBit ? 1'h0 : _GEN_1457; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1459 = _GEN_6085 == 10'h269 ? _GEN_1458 : _GEN_1457; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1460 = io_inputBit | _GEN_1459; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1461 = _GEN_6085 == 10'h269 ? _GEN_1460 : _GEN_1459; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1462 = ~io_inputBit | _GEN_1461; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1463 = _GEN_6085 == 10'h26b ? _GEN_1462 : _GEN_1461; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1464 = io_inputBit ? 1'h0 : _GEN_1463; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1465 = _GEN_6085 == 10'h26b ? _GEN_1464 : _GEN_1463; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1466 = ~io_inputBit ? 1'h0 : _GEN_1465; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1467 = _GEN_6085 == 10'h26d ? _GEN_1466 : _GEN_1465; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1468 = io_inputBit | _GEN_1467; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1469 = _GEN_6085 == 10'h26d ? _GEN_1468 : _GEN_1467; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1470 = ~io_inputBit | _GEN_1469; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1471 = _GEN_6085 == 10'h26f ? _GEN_1470 : _GEN_1469; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1472 = io_inputBit ? 1'h0 : _GEN_1471; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1473 = _GEN_6085 == 10'h26f ? _GEN_1472 : _GEN_1471; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1474 = ~io_inputBit ? 1'h0 : _GEN_1473; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1475 = _GEN_6085 == 10'h271 ? _GEN_1474 : _GEN_1473; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1476 = io_inputBit | _GEN_1475; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1477 = _GEN_6085 == 10'h271 ? _GEN_1476 : _GEN_1475; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1478 = ~io_inputBit | _GEN_1477; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1479 = _GEN_6085 == 10'h273 ? _GEN_1478 : _GEN_1477; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1480 = io_inputBit ? 1'h0 : _GEN_1479; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1481 = _GEN_6085 == 10'h273 ? _GEN_1480 : _GEN_1479; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1482 = ~io_inputBit ? 1'h0 : _GEN_1481; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1483 = _GEN_6085 == 10'h275 ? _GEN_1482 : _GEN_1481; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1484 = io_inputBit | _GEN_1483; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1485 = _GEN_6085 == 10'h275 ? _GEN_1484 : _GEN_1483; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1486 = ~io_inputBit | _GEN_1485; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1487 = _GEN_6085 == 10'h277 ? _GEN_1486 : _GEN_1485; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1488 = io_inputBit ? 1'h0 : _GEN_1487; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1489 = _GEN_6085 == 10'h277 ? _GEN_1488 : _GEN_1487; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1490 = ~io_inputBit ? 1'h0 : _GEN_1489; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1491 = _GEN_6085 == 10'h279 ? _GEN_1490 : _GEN_1489; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1492 = io_inputBit | _GEN_1491; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1493 = _GEN_6085 == 10'h279 ? _GEN_1492 : _GEN_1491; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1494 = ~io_inputBit | _GEN_1493; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1495 = _GEN_6085 == 10'h27b ? _GEN_1494 : _GEN_1493; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1496 = io_inputBit ? 1'h0 : _GEN_1495; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1497 = _GEN_6085 == 10'h27b ? _GEN_1496 : _GEN_1495; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1498 = ~io_inputBit ? 1'h0 : _GEN_1497; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1499 = _GEN_6085 == 10'h27d ? _GEN_1498 : _GEN_1497; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1500 = io_inputBit | _GEN_1499; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1501 = _GEN_6085 == 10'h27d ? _GEN_1500 : _GEN_1499; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1502 = ~io_inputBit | _GEN_1501; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1503 = _GEN_6085 == 10'h27f ? _GEN_1502 : _GEN_1501; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1504 = io_inputBit ? 1'h0 : _GEN_1503; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1505 = _GEN_6085 == 10'h27f ? _GEN_1504 : _GEN_1503; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1506 = ~io_inputBit ? 1'h0 : _GEN_1505; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1507 = _GEN_6085 == 10'h281 ? _GEN_1506 : _GEN_1505; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1508 = io_inputBit | _GEN_1507; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1509 = _GEN_6085 == 10'h281 ? _GEN_1508 : _GEN_1507; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1510 = ~io_inputBit | _GEN_1509; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1511 = _GEN_6085 == 10'h283 ? _GEN_1510 : _GEN_1509; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1512 = io_inputBit ? 1'h0 : _GEN_1511; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1513 = _GEN_6085 == 10'h283 ? _GEN_1512 : _GEN_1511; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1514 = ~io_inputBit ? 1'h0 : _GEN_1513; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1515 = _GEN_6085 == 10'h285 ? _GEN_1514 : _GEN_1513; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1516 = io_inputBit | _GEN_1515; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1517 = _GEN_6085 == 10'h285 ? _GEN_1516 : _GEN_1515; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1518 = ~io_inputBit | _GEN_1517; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1519 = _GEN_6085 == 10'h287 ? _GEN_1518 : _GEN_1517; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1520 = io_inputBit ? 1'h0 : _GEN_1519; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1521 = _GEN_6085 == 10'h287 ? _GEN_1520 : _GEN_1519; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1522 = ~io_inputBit ? 1'h0 : _GEN_1521; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1523 = _GEN_6085 == 10'h289 ? _GEN_1522 : _GEN_1521; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1524 = io_inputBit | _GEN_1523; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1525 = _GEN_6085 == 10'h289 ? _GEN_1524 : _GEN_1523; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1526 = ~io_inputBit | _GEN_1525; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1527 = _GEN_6085 == 10'h28b ? _GEN_1526 : _GEN_1525; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1528 = io_inputBit ? 1'h0 : _GEN_1527; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1529 = _GEN_6085 == 10'h28b ? _GEN_1528 : _GEN_1527; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1530 = ~io_inputBit ? 1'h0 : _GEN_1529; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1531 = _GEN_6085 == 10'h28d ? _GEN_1530 : _GEN_1529; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1532 = io_inputBit | _GEN_1531; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1533 = _GEN_6085 == 10'h28d ? _GEN_1532 : _GEN_1531; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1534 = ~io_inputBit | _GEN_1533; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1535 = _GEN_6085 == 10'h28f ? _GEN_1534 : _GEN_1533; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1536 = io_inputBit ? 1'h0 : _GEN_1535; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1537 = _GEN_6085 == 10'h28f ? _GEN_1536 : _GEN_1535; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1538 = ~io_inputBit ? 1'h0 : _GEN_1537; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1539 = _GEN_6085 == 10'h291 ? _GEN_1538 : _GEN_1537; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1540 = io_inputBit | _GEN_1539; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1541 = _GEN_6085 == 10'h291 ? _GEN_1540 : _GEN_1539; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1542 = ~io_inputBit | _GEN_1541; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1543 = _GEN_6085 == 10'h293 ? _GEN_1542 : _GEN_1541; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1544 = io_inputBit ? 1'h0 : _GEN_1543; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1545 = _GEN_6085 == 10'h293 ? _GEN_1544 : _GEN_1543; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1546 = io_inputBit ? 1'h0 : _GEN_633; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1547 = i == 8'h0 ? _GEN_1546 : _GEN_633; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1548 = io_inputBit ? 1'h0 : _GEN_1547; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1549 = i == 8'h4 ? _GEN_1548 : _GEN_1547; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1550 = io_inputBit ? 1'h0 : _GEN_1549; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1551 = i == 8'h9 ? _GEN_1550 : _GEN_1549; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1552 = ~io_inputBit ? 1'h0 : _GEN_1551; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1553 = i == 8'hf ? _GEN_1552 : _GEN_1551; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1554 = io_inputBit ? 1'h0 : _GEN_1553; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1555 = i == 8'h11 ? _GEN_1554 : _GEN_1553; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1556 = ~io_inputBit ? 1'h0 : _GEN_1555; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1557 = i == 8'h20 ? _GEN_1556 : _GEN_1555; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1558 = io_inputBit ? 1'h0 : _GEN_1557; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1559 = i == 8'h28 ? _GEN_1558 : _GEN_1557; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1560 = io_inputBit ? 1'h0 : _GEN_1559; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1561 = i == 8'h48 ? _GEN_1560 : _GEN_1559; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1562 = ~io_inputBit ? 1'h0 : _GEN_1561; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1563 = i == 8'h4b ? _GEN_1562 : _GEN_1561; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1564 = ~io_inputBit ? 1'h0 : _GEN_1563; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1565 = i == 8'h85 ? _GEN_1564 : _GEN_1563; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1566 = io_inputBit ? 1'h0 : _GEN_1565; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1567 = i == 8'ha4 ? _GEN_1566 : _GEN_1565; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1568 = ~io_inputBit | _GEN_1567; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1569 = _GEN_6084 == 9'h10c ? _GEN_1568 : _GEN_1567; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1570 = io_inputBit ? 1'h0 : _GEN_1569; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1571 = _GEN_6084 == 9'h10c ? _GEN_1570 : _GEN_1569; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1572 = ~io_inputBit | _GEN_1571; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1573 = _GEN_6084 == 9'h10d ? _GEN_1572 : _GEN_1571; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1574 = io_inputBit ? 1'h0 : _GEN_1573; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1575 = _GEN_6084 == 9'h10d ? _GEN_1574 : _GEN_1573; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1576 = ~io_inputBit | _GEN_1575; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1577 = _GEN_6084 == 9'h10e ? _GEN_1576 : _GEN_1575; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1578 = io_inputBit ? 1'h0 : _GEN_1577; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1579 = _GEN_6084 == 9'h10e ? _GEN_1578 : _GEN_1577; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1580 = ~io_inputBit | _GEN_1579; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1581 = _GEN_6084 == 9'h10f ? _GEN_1580 : _GEN_1579; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1582 = io_inputBit ? 1'h0 : _GEN_1581; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1583 = _GEN_6084 == 9'h10f ? _GEN_1582 : _GEN_1581; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1584 = ~io_inputBit | _GEN_1583; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1585 = _GEN_6084 == 9'h110 ? _GEN_1584 : _GEN_1583; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1586 = io_inputBit ? 1'h0 : _GEN_1585; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1587 = _GEN_6084 == 9'h110 ? _GEN_1586 : _GEN_1585; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1588 = ~io_inputBit | _GEN_1587; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1589 = _GEN_6084 == 9'h111 ? _GEN_1588 : _GEN_1587; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1590 = io_inputBit ? 1'h0 : _GEN_1589; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1591 = _GEN_6084 == 9'h111 ? _GEN_1590 : _GEN_1589; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1592 = ~io_inputBit | _GEN_1591; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1593 = _GEN_6084 == 9'h112 ? _GEN_1592 : _GEN_1591; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1594 = io_inputBit ? 1'h0 : _GEN_1593; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1595 = _GEN_6084 == 9'h112 ? _GEN_1594 : _GEN_1593; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1596 = ~io_inputBit | _GEN_1595; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1597 = _GEN_6084 == 9'h113 ? _GEN_1596 : _GEN_1595; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1598 = io_inputBit ? 1'h0 : _GEN_1597; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1599 = _GEN_6084 == 9'h113 ? _GEN_1598 : _GEN_1597; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1600 = ~io_inputBit | _GEN_1599; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1601 = _GEN_6084 == 9'h114 ? _GEN_1600 : _GEN_1599; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1602 = io_inputBit ? 1'h0 : _GEN_1601; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1603 = _GEN_6084 == 9'h114 ? _GEN_1602 : _GEN_1601; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1604 = ~io_inputBit | _GEN_1603; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1605 = _GEN_6084 == 9'h115 ? _GEN_1604 : _GEN_1603; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1606 = io_inputBit ? 1'h0 : _GEN_1605; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1607 = _GEN_6084 == 9'h115 ? _GEN_1606 : _GEN_1605; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1608 = ~io_inputBit | _GEN_1607; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1609 = _GEN_6084 == 9'h116 ? _GEN_1608 : _GEN_1607; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1610 = io_inputBit ? 1'h0 : _GEN_1609; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1611 = _GEN_6084 == 9'h116 ? _GEN_1610 : _GEN_1609; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1612 = ~io_inputBit | _GEN_1611; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1613 = _GEN_6084 == 9'h117 ? _GEN_1612 : _GEN_1611; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1614 = io_inputBit ? 1'h0 : _GEN_1613; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1615 = _GEN_6084 == 9'h117 ? _GEN_1614 : _GEN_1613; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1616 = ~io_inputBit | _GEN_1615; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1617 = _GEN_6084 == 9'h118 ? _GEN_1616 : _GEN_1615; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1618 = io_inputBit ? 1'h0 : _GEN_1617; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1619 = _GEN_6084 == 9'h118 ? _GEN_1618 : _GEN_1617; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1620 = ~io_inputBit | _GEN_1619; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1621 = _GEN_6084 == 9'h119 ? _GEN_1620 : _GEN_1619; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1622 = io_inputBit ? 1'h0 : _GEN_1621; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1623 = _GEN_6084 == 9'h119 ? _GEN_1622 : _GEN_1621; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1624 = ~io_inputBit | _GEN_1623; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1625 = _GEN_6084 == 9'h11a ? _GEN_1624 : _GEN_1623; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1626 = io_inputBit ? 1'h0 : _GEN_1625; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1627 = _GEN_6084 == 9'h11a ? _GEN_1626 : _GEN_1625; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1628 = ~io_inputBit | _GEN_1627; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1629 = _GEN_6084 == 9'h11b ? _GEN_1628 : _GEN_1627; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1630 = io_inputBit ? 1'h0 : _GEN_1629; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1631 = _GEN_6084 == 9'h11b ? _GEN_1630 : _GEN_1629; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1632 = ~io_inputBit | _GEN_1631; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1633 = _GEN_6084 == 9'h11c ? _GEN_1632 : _GEN_1631; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1634 = io_inputBit ? 1'h0 : _GEN_1633; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1635 = _GEN_6084 == 9'h11c ? _GEN_1634 : _GEN_1633; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1636 = ~io_inputBit | _GEN_1635; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1637 = _GEN_6084 == 9'h11d ? _GEN_1636 : _GEN_1635; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1638 = io_inputBit ? 1'h0 : _GEN_1637; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1639 = _GEN_6084 == 9'h11d ? _GEN_1638 : _GEN_1637; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1640 = ~io_inputBit | _GEN_1639; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1641 = _GEN_6084 == 9'h11e ? _GEN_1640 : _GEN_1639; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1642 = io_inputBit ? 1'h0 : _GEN_1641; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1643 = _GEN_6084 == 9'h11e ? _GEN_1642 : _GEN_1641; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1644 = ~io_inputBit | _GEN_1643; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1645 = _GEN_6084 == 9'h11f ? _GEN_1644 : _GEN_1643; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1646 = io_inputBit ? 1'h0 : _GEN_1645; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1647 = _GEN_6084 == 9'h11f ? _GEN_1646 : _GEN_1645; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1648 = ~io_inputBit | _GEN_1647; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1649 = _GEN_6084 == 9'h120 ? _GEN_1648 : _GEN_1647; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1650 = io_inputBit ? 1'h0 : _GEN_1649; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1651 = _GEN_6084 == 9'h120 ? _GEN_1650 : _GEN_1649; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1652 = ~io_inputBit | _GEN_1651; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1653 = _GEN_6084 == 9'h121 ? _GEN_1652 : _GEN_1651; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1654 = io_inputBit ? 1'h0 : _GEN_1653; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1655 = _GEN_6084 == 9'h121 ? _GEN_1654 : _GEN_1653; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1656 = ~io_inputBit | _GEN_1655; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1657 = _GEN_6084 == 9'h122 ? _GEN_1656 : _GEN_1655; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1658 = io_inputBit ? 1'h0 : _GEN_1657; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1659 = _GEN_6084 == 9'h122 ? _GEN_1658 : _GEN_1657; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1660 = ~io_inputBit | _GEN_1659; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1661 = _GEN_6084 == 9'h123 ? _GEN_1660 : _GEN_1659; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1662 = io_inputBit ? 1'h0 : _GEN_1661; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1663 = _GEN_6084 == 9'h123 ? _GEN_1662 : _GEN_1661; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1664 = ~io_inputBit | _GEN_1663; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1665 = _GEN_6084 == 9'h124 ? _GEN_1664 : _GEN_1663; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1666 = io_inputBit ? 1'h0 : _GEN_1665; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1667 = _GEN_6084 == 9'h124 ? _GEN_1666 : _GEN_1665; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1668 = ~io_inputBit ? 1'h0 : _GEN_1667; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1669 = _GEN_6085 == 10'h263 ? _GEN_1668 : _GEN_1667; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1670 = io_inputBit | _GEN_1669; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1671 = _GEN_6085 == 10'h263 ? _GEN_1670 : _GEN_1669; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1672 = ~io_inputBit | _GEN_1671; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1673 = _GEN_6085 == 10'h264 ? _GEN_1672 : _GEN_1671; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1674 = io_inputBit ? 1'h0 : _GEN_1673; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1675 = _GEN_6085 == 10'h264 ? _GEN_1674 : _GEN_1673; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1676 = ~io_inputBit ? 1'h0 : _GEN_1675; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1677 = _GEN_6085 == 10'h265 ? _GEN_1676 : _GEN_1675; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1678 = io_inputBit | _GEN_1677; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1679 = _GEN_6085 == 10'h265 ? _GEN_1678 : _GEN_1677; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1680 = ~io_inputBit | _GEN_1679; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1681 = _GEN_6085 == 10'h266 ? _GEN_1680 : _GEN_1679; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1682 = io_inputBit ? 1'h0 : _GEN_1681; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1683 = _GEN_6085 == 10'h266 ? _GEN_1682 : _GEN_1681; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1684 = ~io_inputBit ? 1'h0 : _GEN_1683; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1685 = _GEN_6085 == 10'h267 ? _GEN_1684 : _GEN_1683; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1686 = io_inputBit | _GEN_1685; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1687 = _GEN_6085 == 10'h267 ? _GEN_1686 : _GEN_1685; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1688 = ~io_inputBit | _GEN_1687; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1689 = _GEN_6085 == 10'h268 ? _GEN_1688 : _GEN_1687; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1690 = io_inputBit ? 1'h0 : _GEN_1689; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1691 = _GEN_6085 == 10'h268 ? _GEN_1690 : _GEN_1689; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1692 = ~io_inputBit ? 1'h0 : _GEN_1691; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1693 = _GEN_6085 == 10'h269 ? _GEN_1692 : _GEN_1691; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1694 = io_inputBit | _GEN_1693; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1695 = _GEN_6085 == 10'h269 ? _GEN_1694 : _GEN_1693; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1696 = ~io_inputBit | _GEN_1695; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1697 = _GEN_6085 == 10'h26a ? _GEN_1696 : _GEN_1695; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1698 = io_inputBit ? 1'h0 : _GEN_1697; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1699 = _GEN_6085 == 10'h26a ? _GEN_1698 : _GEN_1697; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1700 = ~io_inputBit ? 1'h0 : _GEN_1699; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1701 = _GEN_6085 == 10'h26b ? _GEN_1700 : _GEN_1699; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1702 = io_inputBit | _GEN_1701; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1703 = _GEN_6085 == 10'h26b ? _GEN_1702 : _GEN_1701; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1704 = ~io_inputBit | _GEN_1703; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1705 = _GEN_6085 == 10'h26c ? _GEN_1704 : _GEN_1703; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1706 = io_inputBit ? 1'h0 : _GEN_1705; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1707 = _GEN_6085 == 10'h26c ? _GEN_1706 : _GEN_1705; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1708 = ~io_inputBit ? 1'h0 : _GEN_1707; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1709 = _GEN_6085 == 10'h26d ? _GEN_1708 : _GEN_1707; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1710 = io_inputBit | _GEN_1709; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1711 = _GEN_6085 == 10'h26d ? _GEN_1710 : _GEN_1709; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1712 = ~io_inputBit | _GEN_1711; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1713 = _GEN_6085 == 10'h26e ? _GEN_1712 : _GEN_1711; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1714 = io_inputBit ? 1'h0 : _GEN_1713; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1715 = _GEN_6085 == 10'h26e ? _GEN_1714 : _GEN_1713; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1716 = ~io_inputBit ? 1'h0 : _GEN_1715; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1717 = _GEN_6085 == 10'h26f ? _GEN_1716 : _GEN_1715; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1718 = io_inputBit | _GEN_1717; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1719 = _GEN_6085 == 10'h26f ? _GEN_1718 : _GEN_1717; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1720 = ~io_inputBit | _GEN_1719; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1721 = _GEN_6085 == 10'h270 ? _GEN_1720 : _GEN_1719; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1722 = io_inputBit ? 1'h0 : _GEN_1721; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1723 = _GEN_6085 == 10'h270 ? _GEN_1722 : _GEN_1721; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1724 = ~io_inputBit ? 1'h0 : _GEN_1723; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1725 = _GEN_6085 == 10'h271 ? _GEN_1724 : _GEN_1723; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1726 = io_inputBit | _GEN_1725; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1727 = _GEN_6085 == 10'h271 ? _GEN_1726 : _GEN_1725; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1728 = ~io_inputBit | _GEN_1727; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1729 = _GEN_6085 == 10'h272 ? _GEN_1728 : _GEN_1727; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1730 = io_inputBit ? 1'h0 : _GEN_1729; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1731 = _GEN_6085 == 10'h272 ? _GEN_1730 : _GEN_1729; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1732 = ~io_inputBit ? 1'h0 : _GEN_1731; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1733 = _GEN_6085 == 10'h273 ? _GEN_1732 : _GEN_1731; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1734 = io_inputBit | _GEN_1733; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1735 = _GEN_6085 == 10'h273 ? _GEN_1734 : _GEN_1733; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1736 = ~io_inputBit | _GEN_1735; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1737 = _GEN_6085 == 10'h274 ? _GEN_1736 : _GEN_1735; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1738 = io_inputBit ? 1'h0 : _GEN_1737; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1739 = _GEN_6085 == 10'h274 ? _GEN_1738 : _GEN_1737; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1740 = ~io_inputBit ? 1'h0 : _GEN_1739; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1741 = _GEN_6085 == 10'h275 ? _GEN_1740 : _GEN_1739; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1742 = io_inputBit | _GEN_1741; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1743 = _GEN_6085 == 10'h275 ? _GEN_1742 : _GEN_1741; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1744 = ~io_inputBit | _GEN_1743; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1745 = _GEN_6085 == 10'h276 ? _GEN_1744 : _GEN_1743; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1746 = io_inputBit ? 1'h0 : _GEN_1745; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1747 = _GEN_6085 == 10'h276 ? _GEN_1746 : _GEN_1745; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1748 = ~io_inputBit ? 1'h0 : _GEN_1747; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1749 = _GEN_6085 == 10'h277 ? _GEN_1748 : _GEN_1747; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1750 = io_inputBit | _GEN_1749; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1751 = _GEN_6085 == 10'h277 ? _GEN_1750 : _GEN_1749; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1752 = ~io_inputBit | _GEN_1751; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1753 = _GEN_6085 == 10'h278 ? _GEN_1752 : _GEN_1751; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1754 = io_inputBit ? 1'h0 : _GEN_1753; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1755 = _GEN_6085 == 10'h278 ? _GEN_1754 : _GEN_1753; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1756 = ~io_inputBit ? 1'h0 : _GEN_1755; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1757 = _GEN_6085 == 10'h279 ? _GEN_1756 : _GEN_1755; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1758 = io_inputBit | _GEN_1757; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1759 = _GEN_6085 == 10'h279 ? _GEN_1758 : _GEN_1757; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1760 = ~io_inputBit | _GEN_1759; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1761 = _GEN_6085 == 10'h27a ? _GEN_1760 : _GEN_1759; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1762 = io_inputBit ? 1'h0 : _GEN_1761; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1763 = _GEN_6085 == 10'h27a ? _GEN_1762 : _GEN_1761; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1764 = ~io_inputBit ? 1'h0 : _GEN_1763; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1765 = _GEN_6085 == 10'h27b ? _GEN_1764 : _GEN_1763; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1766 = io_inputBit | _GEN_1765; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1767 = _GEN_6085 == 10'h27b ? _GEN_1766 : _GEN_1765; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1768 = ~io_inputBit | _GEN_1767; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1769 = _GEN_6085 == 10'h27c ? _GEN_1768 : _GEN_1767; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1770 = io_inputBit ? 1'h0 : _GEN_1769; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1771 = _GEN_6085 == 10'h27c ? _GEN_1770 : _GEN_1769; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1772 = ~io_inputBit ? 1'h0 : _GEN_1771; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1773 = _GEN_6085 == 10'h27d ? _GEN_1772 : _GEN_1771; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1774 = io_inputBit | _GEN_1773; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1775 = _GEN_6085 == 10'h27d ? _GEN_1774 : _GEN_1773; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1776 = ~io_inputBit | _GEN_1775; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1777 = _GEN_6085 == 10'h27e ? _GEN_1776 : _GEN_1775; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1778 = io_inputBit ? 1'h0 : _GEN_1777; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1779 = _GEN_6085 == 10'h27e ? _GEN_1778 : _GEN_1777; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1780 = ~io_inputBit ? 1'h0 : _GEN_1779; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1781 = _GEN_6085 == 10'h27f ? _GEN_1780 : _GEN_1779; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1782 = io_inputBit | _GEN_1781; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1783 = _GEN_6085 == 10'h27f ? _GEN_1782 : _GEN_1781; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1784 = ~io_inputBit | _GEN_1783; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1785 = _GEN_6085 == 10'h280 ? _GEN_1784 : _GEN_1783; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1786 = io_inputBit ? 1'h0 : _GEN_1785; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1787 = _GEN_6085 == 10'h280 ? _GEN_1786 : _GEN_1785; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1788 = ~io_inputBit ? 1'h0 : _GEN_1787; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1789 = _GEN_6085 == 10'h281 ? _GEN_1788 : _GEN_1787; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1790 = io_inputBit | _GEN_1789; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1791 = _GEN_6085 == 10'h281 ? _GEN_1790 : _GEN_1789; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1792 = ~io_inputBit | _GEN_1791; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1793 = _GEN_6085 == 10'h282 ? _GEN_1792 : _GEN_1791; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1794 = io_inputBit ? 1'h0 : _GEN_1793; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1795 = _GEN_6085 == 10'h282 ? _GEN_1794 : _GEN_1793; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1796 = ~io_inputBit ? 1'h0 : _GEN_1795; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1797 = _GEN_6085 == 10'h283 ? _GEN_1796 : _GEN_1795; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1798 = io_inputBit | _GEN_1797; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1799 = _GEN_6085 == 10'h283 ? _GEN_1798 : _GEN_1797; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1800 = ~io_inputBit | _GEN_1799; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1801 = _GEN_6085 == 10'h284 ? _GEN_1800 : _GEN_1799; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1802 = io_inputBit ? 1'h0 : _GEN_1801; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1803 = _GEN_6085 == 10'h284 ? _GEN_1802 : _GEN_1801; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1804 = ~io_inputBit ? 1'h0 : _GEN_1803; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1805 = _GEN_6085 == 10'h285 ? _GEN_1804 : _GEN_1803; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1806 = io_inputBit | _GEN_1805; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1807 = _GEN_6085 == 10'h285 ? _GEN_1806 : _GEN_1805; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1808 = ~io_inputBit | _GEN_1807; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1809 = _GEN_6085 == 10'h286 ? _GEN_1808 : _GEN_1807; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1810 = io_inputBit ? 1'h0 : _GEN_1809; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1811 = _GEN_6085 == 10'h286 ? _GEN_1810 : _GEN_1809; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1812 = ~io_inputBit ? 1'h0 : _GEN_1811; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1813 = _GEN_6085 == 10'h287 ? _GEN_1812 : _GEN_1811; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1814 = io_inputBit | _GEN_1813; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1815 = _GEN_6085 == 10'h287 ? _GEN_1814 : _GEN_1813; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1816 = ~io_inputBit | _GEN_1815; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1817 = _GEN_6085 == 10'h288 ? _GEN_1816 : _GEN_1815; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1818 = io_inputBit ? 1'h0 : _GEN_1817; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1819 = _GEN_6085 == 10'h288 ? _GEN_1818 : _GEN_1817; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1820 = ~io_inputBit ? 1'h0 : _GEN_1819; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1821 = _GEN_6085 == 10'h289 ? _GEN_1820 : _GEN_1819; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1822 = io_inputBit | _GEN_1821; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1823 = _GEN_6085 == 10'h289 ? _GEN_1822 : _GEN_1821; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1824 = ~io_inputBit | _GEN_1823; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1825 = _GEN_6085 == 10'h28a ? _GEN_1824 : _GEN_1823; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1826 = io_inputBit ? 1'h0 : _GEN_1825; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1827 = _GEN_6085 == 10'h28a ? _GEN_1826 : _GEN_1825; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1828 = ~io_inputBit ? 1'h0 : _GEN_1827; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1829 = _GEN_6085 == 10'h28b ? _GEN_1828 : _GEN_1827; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1830 = io_inputBit | _GEN_1829; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1831 = _GEN_6085 == 10'h28b ? _GEN_1830 : _GEN_1829; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1832 = ~io_inputBit | _GEN_1831; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1833 = _GEN_6085 == 10'h28c ? _GEN_1832 : _GEN_1831; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1834 = io_inputBit ? 1'h0 : _GEN_1833; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1835 = _GEN_6085 == 10'h28c ? _GEN_1834 : _GEN_1833; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1836 = ~io_inputBit ? 1'h0 : _GEN_1835; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1837 = _GEN_6085 == 10'h28d ? _GEN_1836 : _GEN_1835; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1838 = io_inputBit | _GEN_1837; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1839 = _GEN_6085 == 10'h28d ? _GEN_1838 : _GEN_1837; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1840 = ~io_inputBit | _GEN_1839; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1841 = _GEN_6085 == 10'h28e ? _GEN_1840 : _GEN_1839; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1842 = io_inputBit ? 1'h0 : _GEN_1841; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1843 = _GEN_6085 == 10'h28e ? _GEN_1842 : _GEN_1841; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1844 = ~io_inputBit ? 1'h0 : _GEN_1843; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1845 = _GEN_6085 == 10'h28f ? _GEN_1844 : _GEN_1843; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1846 = io_inputBit | _GEN_1845; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1847 = _GEN_6085 == 10'h28f ? _GEN_1846 : _GEN_1845; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1848 = ~io_inputBit | _GEN_1847; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1849 = _GEN_6085 == 10'h290 ? _GEN_1848 : _GEN_1847; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1850 = io_inputBit ? 1'h0 : _GEN_1849; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1851 = _GEN_6085 == 10'h290 ? _GEN_1850 : _GEN_1849; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1852 = ~io_inputBit ? 1'h0 : _GEN_1851; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1853 = _GEN_6085 == 10'h291 ? _GEN_1852 : _GEN_1851; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1854 = io_inputBit | _GEN_1853; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1855 = _GEN_6085 == 10'h291 ? _GEN_1854 : _GEN_1853; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1856 = ~io_inputBit | _GEN_1855; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1857 = _GEN_6085 == 10'h292 ? _GEN_1856 : _GEN_1855; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1858 = io_inputBit ? 1'h0 : _GEN_1857; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1859 = _GEN_6085 == 10'h292 ? _GEN_1858 : _GEN_1857; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1860 = ~io_inputBit ? 1'h0 : _GEN_1859; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1861 = _GEN_6085 == 10'h293 ? _GEN_1860 : _GEN_1859; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1862 = io_inputBit | _GEN_1861; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1863 = _GEN_6085 == 10'h293 ? _GEN_1862 : _GEN_1861; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1864 = ~io_inputBit | _GEN_1863; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1865 = _GEN_6085 == 10'h294 ? _GEN_1864 : _GEN_1863; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1866 = io_inputBit ? 1'h0 : _GEN_1865; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1867 = _GEN_6085 == 10'h294 ? _GEN_1866 : _GEN_1865; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1868 = io_inputBit ? 1'h0 : _GEN_851; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1869 = i == 8'h0 ? _GEN_1868 : _GEN_851; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1870 = io_inputBit ? 1'h0 : _GEN_1869; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1871 = i == 8'h4 ? _GEN_1870 : _GEN_1869; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1872 = io_inputBit ? 1'h0 : _GEN_1871; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1873 = i == 8'h9 ? _GEN_1872 : _GEN_1871; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1874 = ~io_inputBit ? 1'h0 : _GEN_1873; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1875 = i == 8'hf ? _GEN_1874 : _GEN_1873; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1876 = io_inputBit ? 1'h0 : _GEN_1875; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1877 = i == 8'h11 ? _GEN_1876 : _GEN_1875; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1878 = ~io_inputBit ? 1'h0 : _GEN_1877; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1879 = i == 8'h20 ? _GEN_1878 : _GEN_1877; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1880 = io_inputBit ? 1'h0 : _GEN_1879; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1881 = i == 8'h28 ? _GEN_1880 : _GEN_1879; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1882 = io_inputBit ? 1'h0 : _GEN_1881; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1883 = i == 8'h48 ? _GEN_1882 : _GEN_1881; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1884 = ~io_inputBit ? 1'h0 : _GEN_1883; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1885 = i == 8'h4b ? _GEN_1884 : _GEN_1883; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1886 = io_inputBit ? 1'h0 : _GEN_1885; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1887 = i == 8'ha4 ? _GEN_1886 : _GEN_1885; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1888 = ~io_inputBit ? 1'h0 : _GEN_1887; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1889 = _GEN_6084 == 9'h10b ? _GEN_1888 : _GEN_1887; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1890 = io_inputBit ? 1'h0 : _GEN_1889; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1891 = _GEN_6084 == 9'h124 ? _GEN_1890 : _GEN_1889; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1892 = ~io_inputBit ? 1'h0 : _GEN_1891; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1893 = _GEN_6085 == 10'h218 ? _GEN_1892 : _GEN_1891; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1894 = io_inputBit | _GEN_1893; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1895 = _GEN_6085 == 10'h218 ? _GEN_1894 : _GEN_1893; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1896 = ~io_inputBit ? 1'h0 : _GEN_1895; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1897 = _GEN_6085 == 10'h219 ? _GEN_1896 : _GEN_1895; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1898 = io_inputBit | _GEN_1897; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1899 = _GEN_6085 == 10'h219 ? _GEN_1898 : _GEN_1897; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1900 = ~io_inputBit ? 1'h0 : _GEN_1899; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1901 = _GEN_6085 == 10'h21a ? _GEN_1900 : _GEN_1899; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1902 = io_inputBit | _GEN_1901; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1903 = _GEN_6085 == 10'h21a ? _GEN_1902 : _GEN_1901; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1904 = ~io_inputBit ? 1'h0 : _GEN_1903; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1905 = _GEN_6085 == 10'h21b ? _GEN_1904 : _GEN_1903; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1906 = io_inputBit | _GEN_1905; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1907 = _GEN_6085 == 10'h21b ? _GEN_1906 : _GEN_1905; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1908 = ~io_inputBit ? 1'h0 : _GEN_1907; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1909 = _GEN_6085 == 10'h21c ? _GEN_1908 : _GEN_1907; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1910 = io_inputBit | _GEN_1909; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1911 = _GEN_6085 == 10'h21c ? _GEN_1910 : _GEN_1909; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1912 = ~io_inputBit ? 1'h0 : _GEN_1911; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1913 = _GEN_6085 == 10'h21d ? _GEN_1912 : _GEN_1911; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1914 = io_inputBit | _GEN_1913; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1915 = _GEN_6085 == 10'h21d ? _GEN_1914 : _GEN_1913; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1916 = ~io_inputBit ? 1'h0 : _GEN_1915; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1917 = _GEN_6085 == 10'h21e ? _GEN_1916 : _GEN_1915; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1918 = io_inputBit | _GEN_1917; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1919 = _GEN_6085 == 10'h21e ? _GEN_1918 : _GEN_1917; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1920 = ~io_inputBit ? 1'h0 : _GEN_1919; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1921 = _GEN_6085 == 10'h21f ? _GEN_1920 : _GEN_1919; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1922 = io_inputBit | _GEN_1921; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1923 = _GEN_6085 == 10'h21f ? _GEN_1922 : _GEN_1921; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1924 = ~io_inputBit ? 1'h0 : _GEN_1923; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1925 = _GEN_6085 == 10'h220 ? _GEN_1924 : _GEN_1923; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1926 = io_inputBit | _GEN_1925; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1927 = _GEN_6085 == 10'h220 ? _GEN_1926 : _GEN_1925; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1928 = ~io_inputBit ? 1'h0 : _GEN_1927; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1929 = _GEN_6085 == 10'h221 ? _GEN_1928 : _GEN_1927; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1930 = io_inputBit | _GEN_1929; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1931 = _GEN_6085 == 10'h221 ? _GEN_1930 : _GEN_1929; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1932 = ~io_inputBit ? 1'h0 : _GEN_1931; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1933 = _GEN_6085 == 10'h222 ? _GEN_1932 : _GEN_1931; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1934 = io_inputBit | _GEN_1933; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1935 = _GEN_6085 == 10'h222 ? _GEN_1934 : _GEN_1933; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1936 = ~io_inputBit ? 1'h0 : _GEN_1935; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1937 = _GEN_6085 == 10'h223 ? _GEN_1936 : _GEN_1935; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1938 = io_inputBit | _GEN_1937; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1939 = _GEN_6085 == 10'h223 ? _GEN_1938 : _GEN_1937; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1940 = ~io_inputBit ? 1'h0 : _GEN_1939; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1941 = _GEN_6085 == 10'h224 ? _GEN_1940 : _GEN_1939; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1942 = io_inputBit | _GEN_1941; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1943 = _GEN_6085 == 10'h224 ? _GEN_1942 : _GEN_1941; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1944 = ~io_inputBit ? 1'h0 : _GEN_1943; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1945 = _GEN_6085 == 10'h225 ? _GEN_1944 : _GEN_1943; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1946 = io_inputBit | _GEN_1945; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1947 = _GEN_6085 == 10'h225 ? _GEN_1946 : _GEN_1945; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1948 = ~io_inputBit ? 1'h0 : _GEN_1947; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1949 = _GEN_6085 == 10'h226 ? _GEN_1948 : _GEN_1947; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1950 = io_inputBit | _GEN_1949; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1951 = _GEN_6085 == 10'h226 ? _GEN_1950 : _GEN_1949; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1952 = ~io_inputBit ? 1'h0 : _GEN_1951; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1953 = _GEN_6085 == 10'h227 ? _GEN_1952 : _GEN_1951; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1954 = io_inputBit | _GEN_1953; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1955 = _GEN_6085 == 10'h227 ? _GEN_1954 : _GEN_1953; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1956 = ~io_inputBit ? 1'h0 : _GEN_1955; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1957 = _GEN_6085 == 10'h228 ? _GEN_1956 : _GEN_1955; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1958 = io_inputBit | _GEN_1957; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1959 = _GEN_6085 == 10'h228 ? _GEN_1958 : _GEN_1957; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1960 = ~io_inputBit ? 1'h0 : _GEN_1959; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1961 = _GEN_6085 == 10'h229 ? _GEN_1960 : _GEN_1959; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1962 = io_inputBit | _GEN_1961; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1963 = _GEN_6085 == 10'h229 ? _GEN_1962 : _GEN_1961; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1964 = ~io_inputBit ? 1'h0 : _GEN_1963; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1965 = _GEN_6085 == 10'h22a ? _GEN_1964 : _GEN_1963; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1966 = io_inputBit | _GEN_1965; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1967 = _GEN_6085 == 10'h22a ? _GEN_1966 : _GEN_1965; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1968 = ~io_inputBit ? 1'h0 : _GEN_1967; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1969 = _GEN_6085 == 10'h22b ? _GEN_1968 : _GEN_1967; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1970 = io_inputBit | _GEN_1969; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1971 = _GEN_6085 == 10'h22b ? _GEN_1970 : _GEN_1969; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1972 = ~io_inputBit ? 1'h0 : _GEN_1971; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1973 = _GEN_6085 == 10'h22c ? _GEN_1972 : _GEN_1971; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1974 = io_inputBit | _GEN_1973; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1975 = _GEN_6085 == 10'h22c ? _GEN_1974 : _GEN_1973; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1976 = ~io_inputBit ? 1'h0 : _GEN_1975; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1977 = _GEN_6085 == 10'h22d ? _GEN_1976 : _GEN_1975; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1978 = io_inputBit | _GEN_1977; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1979 = _GEN_6085 == 10'h22d ? _GEN_1978 : _GEN_1977; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1980 = ~io_inputBit ? 1'h0 : _GEN_1979; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1981 = _GEN_6085 == 10'h22e ? _GEN_1980 : _GEN_1979; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1982 = io_inputBit | _GEN_1981; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1983 = _GEN_6085 == 10'h22e ? _GEN_1982 : _GEN_1981; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1984 = ~io_inputBit ? 1'h0 : _GEN_1983; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1985 = _GEN_6085 == 10'h22f ? _GEN_1984 : _GEN_1983; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1986 = io_inputBit | _GEN_1985; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1987 = _GEN_6085 == 10'h22f ? _GEN_1986 : _GEN_1985; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1988 = ~io_inputBit ? 1'h0 : _GEN_1987; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1989 = _GEN_6085 == 10'h230 ? _GEN_1988 : _GEN_1987; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1990 = io_inputBit | _GEN_1989; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1991 = _GEN_6085 == 10'h230 ? _GEN_1990 : _GEN_1989; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1992 = ~io_inputBit ? 1'h0 : _GEN_1991; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1993 = _GEN_6085 == 10'h231 ? _GEN_1992 : _GEN_1991; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1994 = io_inputBit | _GEN_1993; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1995 = _GEN_6085 == 10'h231 ? _GEN_1994 : _GEN_1993; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1996 = ~io_inputBit ? 1'h0 : _GEN_1995; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1997 = _GEN_6085 == 10'h232 ? _GEN_1996 : _GEN_1995; // @[lut_mem_online.scala 235:34]
  wire  _GEN_1998 = io_inputBit | _GEN_1997; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_1999 = _GEN_6085 == 10'h232 ? _GEN_1998 : _GEN_1997; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2000 = ~io_inputBit ? 1'h0 : _GEN_1999; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2001 = _GEN_6085 == 10'h233 ? _GEN_2000 : _GEN_1999; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2002 = io_inputBit | _GEN_2001; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2003 = _GEN_6085 == 10'h233 ? _GEN_2002 : _GEN_2001; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2004 = ~io_inputBit ? 1'h0 : _GEN_2003; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2005 = _GEN_6085 == 10'h234 ? _GEN_2004 : _GEN_2003; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2006 = io_inputBit | _GEN_2005; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2007 = _GEN_6085 == 10'h234 ? _GEN_2006 : _GEN_2005; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2008 = ~io_inputBit ? 1'h0 : _GEN_2007; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2009 = _GEN_6085 == 10'h235 ? _GEN_2008 : _GEN_2007; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2010 = io_inputBit | _GEN_2009; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2011 = _GEN_6085 == 10'h235 ? _GEN_2010 : _GEN_2009; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2012 = ~io_inputBit ? 1'h0 : _GEN_2011; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2013 = _GEN_6085 == 10'h236 ? _GEN_2012 : _GEN_2011; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2014 = io_inputBit | _GEN_2013; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2015 = _GEN_6085 == 10'h236 ? _GEN_2014 : _GEN_2013; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2016 = ~io_inputBit ? 1'h0 : _GEN_2015; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2017 = _GEN_6085 == 10'h237 ? _GEN_2016 : _GEN_2015; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2018 = io_inputBit | _GEN_2017; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2019 = _GEN_6085 == 10'h237 ? _GEN_2018 : _GEN_2017; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2020 = ~io_inputBit ? 1'h0 : _GEN_2019; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2021 = _GEN_6085 == 10'h238 ? _GEN_2020 : _GEN_2019; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2022 = io_inputBit | _GEN_2021; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2023 = _GEN_6085 == 10'h238 ? _GEN_2022 : _GEN_2021; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2024 = ~io_inputBit ? 1'h0 : _GEN_2023; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2025 = _GEN_6085 == 10'h239 ? _GEN_2024 : _GEN_2023; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2026 = io_inputBit | _GEN_2025; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2027 = _GEN_6085 == 10'h239 ? _GEN_2026 : _GEN_2025; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2028 = ~io_inputBit ? 1'h0 : _GEN_2027; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2029 = _GEN_6085 == 10'h23a ? _GEN_2028 : _GEN_2027; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2030 = io_inputBit | _GEN_2029; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2031 = _GEN_6085 == 10'h23a ? _GEN_2030 : _GEN_2029; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2032 = ~io_inputBit ? 1'h0 : _GEN_2031; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2033 = _GEN_6085 == 10'h23b ? _GEN_2032 : _GEN_2031; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2034 = io_inputBit | _GEN_2033; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2035 = _GEN_6085 == 10'h23b ? _GEN_2034 : _GEN_2033; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2036 = ~io_inputBit ? 1'h0 : _GEN_2035; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2037 = _GEN_6085 == 10'h23c ? _GEN_2036 : _GEN_2035; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2038 = io_inputBit | _GEN_2037; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2039 = _GEN_6085 == 10'h23c ? _GEN_2038 : _GEN_2037; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2040 = ~io_inputBit ? 1'h0 : _GEN_2039; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2041 = _GEN_6085 == 10'h23d ? _GEN_2040 : _GEN_2039; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2042 = io_inputBit | _GEN_2041; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2043 = _GEN_6085 == 10'h23d ? _GEN_2042 : _GEN_2041; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2044 = ~io_inputBit ? 1'h0 : _GEN_2043; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2045 = _GEN_6085 == 10'h23e ? _GEN_2044 : _GEN_2043; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2046 = io_inputBit | _GEN_2045; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2047 = _GEN_6085 == 10'h23e ? _GEN_2046 : _GEN_2045; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2048 = ~io_inputBit ? 1'h0 : _GEN_2047; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2049 = _GEN_6085 == 10'h23f ? _GEN_2048 : _GEN_2047; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2050 = io_inputBit | _GEN_2049; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2051 = _GEN_6085 == 10'h23f ? _GEN_2050 : _GEN_2049; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2052 = ~io_inputBit ? 1'h0 : _GEN_2051; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2053 = _GEN_6085 == 10'h240 ? _GEN_2052 : _GEN_2051; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2054 = io_inputBit | _GEN_2053; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2055 = _GEN_6085 == 10'h240 ? _GEN_2054 : _GEN_2053; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2056 = ~io_inputBit ? 1'h0 : _GEN_2055; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2057 = _GEN_6085 == 10'h241 ? _GEN_2056 : _GEN_2055; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2058 = io_inputBit | _GEN_2057; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2059 = _GEN_6085 == 10'h241 ? _GEN_2058 : _GEN_2057; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2060 = ~io_inputBit ? 1'h0 : _GEN_2059; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2061 = _GEN_6085 == 10'h242 ? _GEN_2060 : _GEN_2059; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2062 = io_inputBit | _GEN_2061; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2063 = _GEN_6085 == 10'h242 ? _GEN_2062 : _GEN_2061; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2064 = ~io_inputBit ? 1'h0 : _GEN_2063; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2065 = _GEN_6085 == 10'h243 ? _GEN_2064 : _GEN_2063; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2066 = io_inputBit | _GEN_2065; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2067 = _GEN_6085 == 10'h243 ? _GEN_2066 : _GEN_2065; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2068 = ~io_inputBit ? 1'h0 : _GEN_2067; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2069 = _GEN_6085 == 10'h244 ? _GEN_2068 : _GEN_2067; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2070 = io_inputBit | _GEN_2069; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2071 = _GEN_6085 == 10'h244 ? _GEN_2070 : _GEN_2069; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2072 = ~io_inputBit ? 1'h0 : _GEN_2071; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2073 = _GEN_6085 == 10'h245 ? _GEN_2072 : _GEN_2071; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2074 = io_inputBit | _GEN_2073; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2075 = _GEN_6085 == 10'h245 ? _GEN_2074 : _GEN_2073; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2076 = ~io_inputBit ? 1'h0 : _GEN_2075; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2077 = _GEN_6085 == 10'h246 ? _GEN_2076 : _GEN_2075; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2078 = io_inputBit | _GEN_2077; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2079 = _GEN_6085 == 10'h246 ? _GEN_2078 : _GEN_2077; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2080 = ~io_inputBit ? 1'h0 : _GEN_2079; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2081 = _GEN_6085 == 10'h247 ? _GEN_2080 : _GEN_2079; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2082 = io_inputBit | _GEN_2081; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2083 = _GEN_6085 == 10'h247 ? _GEN_2082 : _GEN_2081; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2084 = ~io_inputBit ? 1'h0 : _GEN_2083; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2085 = _GEN_6085 == 10'h248 ? _GEN_2084 : _GEN_2083; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2086 = io_inputBit | _GEN_2085; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2087 = _GEN_6085 == 10'h248 ? _GEN_2086 : _GEN_2085; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2088 = ~io_inputBit ? 1'h0 : _GEN_2087; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2089 = _GEN_6085 == 10'h249 ? _GEN_2088 : _GEN_2087; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2090 = io_inputBit | _GEN_2089; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2091 = _GEN_6085 == 10'h249 ? _GEN_2090 : _GEN_2089; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2092 = ~io_inputBit ? 1'h0 : _GEN_2091; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2093 = _GEN_6085 == 10'h263 ? _GEN_2092 : _GEN_2091; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2094 = io_inputBit | _GEN_2093; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2095 = _GEN_6085 == 10'h263 ? _GEN_2094 : _GEN_2093; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2096 = ~io_inputBit ? 1'h0 : _GEN_2095; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2097 = _GEN_6085 == 10'h264 ? _GEN_2096 : _GEN_2095; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2098 = io_inputBit | _GEN_2097; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2099 = _GEN_6085 == 10'h264 ? _GEN_2098 : _GEN_2097; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2100 = ~io_inputBit ? 1'h0 : _GEN_2099; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2101 = _GEN_6085 == 10'h265 ? _GEN_2100 : _GEN_2099; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2102 = io_inputBit | _GEN_2101; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2103 = _GEN_6085 == 10'h265 ? _GEN_2102 : _GEN_2101; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2104 = ~io_inputBit ? 1'h0 : _GEN_2103; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2105 = _GEN_6085 == 10'h266 ? _GEN_2104 : _GEN_2103; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2106 = io_inputBit | _GEN_2105; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2107 = _GEN_6085 == 10'h266 ? _GEN_2106 : _GEN_2105; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2108 = ~io_inputBit ? 1'h0 : _GEN_2107; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2109 = _GEN_6085 == 10'h267 ? _GEN_2108 : _GEN_2107; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2110 = io_inputBit | _GEN_2109; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2111 = _GEN_6085 == 10'h267 ? _GEN_2110 : _GEN_2109; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2112 = ~io_inputBit ? 1'h0 : _GEN_2111; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2113 = _GEN_6085 == 10'h268 ? _GEN_2112 : _GEN_2111; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2114 = io_inputBit | _GEN_2113; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2115 = _GEN_6085 == 10'h268 ? _GEN_2114 : _GEN_2113; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2116 = ~io_inputBit ? 1'h0 : _GEN_2115; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2117 = _GEN_6085 == 10'h269 ? _GEN_2116 : _GEN_2115; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2118 = io_inputBit | _GEN_2117; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2119 = _GEN_6085 == 10'h269 ? _GEN_2118 : _GEN_2117; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2120 = ~io_inputBit ? 1'h0 : _GEN_2119; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2121 = _GEN_6085 == 10'h26a ? _GEN_2120 : _GEN_2119; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2122 = io_inputBit | _GEN_2121; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2123 = _GEN_6085 == 10'h26a ? _GEN_2122 : _GEN_2121; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2124 = ~io_inputBit ? 1'h0 : _GEN_2123; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2125 = _GEN_6085 == 10'h26b ? _GEN_2124 : _GEN_2123; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2126 = io_inputBit | _GEN_2125; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2127 = _GEN_6085 == 10'h26b ? _GEN_2126 : _GEN_2125; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2128 = ~io_inputBit ? 1'h0 : _GEN_2127; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2129 = _GEN_6085 == 10'h26c ? _GEN_2128 : _GEN_2127; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2130 = io_inputBit | _GEN_2129; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2131 = _GEN_6085 == 10'h26c ? _GEN_2130 : _GEN_2129; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2132 = ~io_inputBit ? 1'h0 : _GEN_2131; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2133 = _GEN_6085 == 10'h26d ? _GEN_2132 : _GEN_2131; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2134 = io_inputBit | _GEN_2133; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2135 = _GEN_6085 == 10'h26d ? _GEN_2134 : _GEN_2133; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2136 = ~io_inputBit ? 1'h0 : _GEN_2135; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2137 = _GEN_6085 == 10'h26e ? _GEN_2136 : _GEN_2135; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2138 = io_inputBit | _GEN_2137; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2139 = _GEN_6085 == 10'h26e ? _GEN_2138 : _GEN_2137; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2140 = ~io_inputBit ? 1'h0 : _GEN_2139; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2141 = _GEN_6085 == 10'h26f ? _GEN_2140 : _GEN_2139; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2142 = io_inputBit | _GEN_2141; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2143 = _GEN_6085 == 10'h26f ? _GEN_2142 : _GEN_2141; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2144 = ~io_inputBit ? 1'h0 : _GEN_2143; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2145 = _GEN_6085 == 10'h270 ? _GEN_2144 : _GEN_2143; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2146 = io_inputBit | _GEN_2145; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2147 = _GEN_6085 == 10'h270 ? _GEN_2146 : _GEN_2145; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2148 = ~io_inputBit ? 1'h0 : _GEN_2147; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2149 = _GEN_6085 == 10'h271 ? _GEN_2148 : _GEN_2147; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2150 = io_inputBit | _GEN_2149; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2151 = _GEN_6085 == 10'h271 ? _GEN_2150 : _GEN_2149; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2152 = ~io_inputBit ? 1'h0 : _GEN_2151; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2153 = _GEN_6085 == 10'h272 ? _GEN_2152 : _GEN_2151; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2154 = io_inputBit | _GEN_2153; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2155 = _GEN_6085 == 10'h272 ? _GEN_2154 : _GEN_2153; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2156 = ~io_inputBit ? 1'h0 : _GEN_2155; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2157 = _GEN_6085 == 10'h273 ? _GEN_2156 : _GEN_2155; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2158 = io_inputBit | _GEN_2157; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2159 = _GEN_6085 == 10'h273 ? _GEN_2158 : _GEN_2157; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2160 = ~io_inputBit ? 1'h0 : _GEN_2159; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2161 = _GEN_6085 == 10'h274 ? _GEN_2160 : _GEN_2159; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2162 = io_inputBit | _GEN_2161; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2163 = _GEN_6085 == 10'h274 ? _GEN_2162 : _GEN_2161; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2164 = ~io_inputBit ? 1'h0 : _GEN_2163; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2165 = _GEN_6085 == 10'h275 ? _GEN_2164 : _GEN_2163; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2166 = io_inputBit | _GEN_2165; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2167 = _GEN_6085 == 10'h275 ? _GEN_2166 : _GEN_2165; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2168 = ~io_inputBit ? 1'h0 : _GEN_2167; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2169 = _GEN_6085 == 10'h276 ? _GEN_2168 : _GEN_2167; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2170 = io_inputBit | _GEN_2169; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2171 = _GEN_6085 == 10'h276 ? _GEN_2170 : _GEN_2169; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2172 = ~io_inputBit ? 1'h0 : _GEN_2171; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2173 = _GEN_6085 == 10'h277 ? _GEN_2172 : _GEN_2171; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2174 = io_inputBit | _GEN_2173; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2175 = _GEN_6085 == 10'h277 ? _GEN_2174 : _GEN_2173; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2176 = ~io_inputBit ? 1'h0 : _GEN_2175; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2177 = _GEN_6085 == 10'h278 ? _GEN_2176 : _GEN_2175; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2178 = io_inputBit | _GEN_2177; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2179 = _GEN_6085 == 10'h278 ? _GEN_2178 : _GEN_2177; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2180 = ~io_inputBit ? 1'h0 : _GEN_2179; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2181 = _GEN_6085 == 10'h279 ? _GEN_2180 : _GEN_2179; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2182 = io_inputBit | _GEN_2181; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2183 = _GEN_6085 == 10'h279 ? _GEN_2182 : _GEN_2181; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2184 = ~io_inputBit ? 1'h0 : _GEN_2183; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2185 = _GEN_6085 == 10'h27a ? _GEN_2184 : _GEN_2183; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2186 = io_inputBit | _GEN_2185; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2187 = _GEN_6085 == 10'h27a ? _GEN_2186 : _GEN_2185; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2188 = ~io_inputBit ? 1'h0 : _GEN_2187; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2189 = _GEN_6085 == 10'h27b ? _GEN_2188 : _GEN_2187; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2190 = io_inputBit | _GEN_2189; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2191 = _GEN_6085 == 10'h27b ? _GEN_2190 : _GEN_2189; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2192 = ~io_inputBit ? 1'h0 : _GEN_2191; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2193 = _GEN_6085 == 10'h27c ? _GEN_2192 : _GEN_2191; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2194 = io_inputBit | _GEN_2193; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2195 = _GEN_6085 == 10'h27c ? _GEN_2194 : _GEN_2193; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2196 = ~io_inputBit ? 1'h0 : _GEN_2195; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2197 = _GEN_6085 == 10'h27d ? _GEN_2196 : _GEN_2195; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2198 = io_inputBit | _GEN_2197; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2199 = _GEN_6085 == 10'h27d ? _GEN_2198 : _GEN_2197; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2200 = ~io_inputBit ? 1'h0 : _GEN_2199; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2201 = _GEN_6085 == 10'h27e ? _GEN_2200 : _GEN_2199; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2202 = io_inputBit | _GEN_2201; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2203 = _GEN_6085 == 10'h27e ? _GEN_2202 : _GEN_2201; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2204 = ~io_inputBit ? 1'h0 : _GEN_2203; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2205 = _GEN_6085 == 10'h27f ? _GEN_2204 : _GEN_2203; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2206 = io_inputBit | _GEN_2205; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2207 = _GEN_6085 == 10'h27f ? _GEN_2206 : _GEN_2205; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2208 = ~io_inputBit ? 1'h0 : _GEN_2207; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2209 = _GEN_6085 == 10'h280 ? _GEN_2208 : _GEN_2207; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2210 = io_inputBit | _GEN_2209; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2211 = _GEN_6085 == 10'h280 ? _GEN_2210 : _GEN_2209; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2212 = ~io_inputBit ? 1'h0 : _GEN_2211; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2213 = _GEN_6085 == 10'h281 ? _GEN_2212 : _GEN_2211; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2214 = io_inputBit | _GEN_2213; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2215 = _GEN_6085 == 10'h281 ? _GEN_2214 : _GEN_2213; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2216 = ~io_inputBit ? 1'h0 : _GEN_2215; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2217 = _GEN_6085 == 10'h282 ? _GEN_2216 : _GEN_2215; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2218 = io_inputBit | _GEN_2217; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2219 = _GEN_6085 == 10'h282 ? _GEN_2218 : _GEN_2217; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2220 = ~io_inputBit ? 1'h0 : _GEN_2219; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2221 = _GEN_6085 == 10'h283 ? _GEN_2220 : _GEN_2219; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2222 = io_inputBit | _GEN_2221; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2223 = _GEN_6085 == 10'h283 ? _GEN_2222 : _GEN_2221; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2224 = ~io_inputBit ? 1'h0 : _GEN_2223; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2225 = _GEN_6085 == 10'h284 ? _GEN_2224 : _GEN_2223; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2226 = io_inputBit | _GEN_2225; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2227 = _GEN_6085 == 10'h284 ? _GEN_2226 : _GEN_2225; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2228 = ~io_inputBit ? 1'h0 : _GEN_2227; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2229 = _GEN_6085 == 10'h285 ? _GEN_2228 : _GEN_2227; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2230 = io_inputBit | _GEN_2229; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2231 = _GEN_6085 == 10'h285 ? _GEN_2230 : _GEN_2229; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2232 = ~io_inputBit ? 1'h0 : _GEN_2231; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2233 = _GEN_6085 == 10'h286 ? _GEN_2232 : _GEN_2231; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2234 = io_inputBit | _GEN_2233; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2235 = _GEN_6085 == 10'h286 ? _GEN_2234 : _GEN_2233; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2236 = ~io_inputBit ? 1'h0 : _GEN_2235; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2237 = _GEN_6085 == 10'h287 ? _GEN_2236 : _GEN_2235; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2238 = io_inputBit | _GEN_2237; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2239 = _GEN_6085 == 10'h287 ? _GEN_2238 : _GEN_2237; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2240 = ~io_inputBit ? 1'h0 : _GEN_2239; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2241 = _GEN_6085 == 10'h288 ? _GEN_2240 : _GEN_2239; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2242 = io_inputBit | _GEN_2241; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2243 = _GEN_6085 == 10'h288 ? _GEN_2242 : _GEN_2241; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2244 = ~io_inputBit ? 1'h0 : _GEN_2243; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2245 = _GEN_6085 == 10'h289 ? _GEN_2244 : _GEN_2243; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2246 = io_inputBit | _GEN_2245; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2247 = _GEN_6085 == 10'h289 ? _GEN_2246 : _GEN_2245; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2248 = ~io_inputBit ? 1'h0 : _GEN_2247; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2249 = _GEN_6085 == 10'h28a ? _GEN_2248 : _GEN_2247; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2250 = io_inputBit | _GEN_2249; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2251 = _GEN_6085 == 10'h28a ? _GEN_2250 : _GEN_2249; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2252 = ~io_inputBit ? 1'h0 : _GEN_2251; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2253 = _GEN_6085 == 10'h28b ? _GEN_2252 : _GEN_2251; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2254 = io_inputBit | _GEN_2253; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2255 = _GEN_6085 == 10'h28b ? _GEN_2254 : _GEN_2253; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2256 = ~io_inputBit ? 1'h0 : _GEN_2255; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2257 = _GEN_6085 == 10'h28c ? _GEN_2256 : _GEN_2255; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2258 = io_inputBit | _GEN_2257; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2259 = _GEN_6085 == 10'h28c ? _GEN_2258 : _GEN_2257; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2260 = ~io_inputBit ? 1'h0 : _GEN_2259; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2261 = _GEN_6085 == 10'h28d ? _GEN_2260 : _GEN_2259; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2262 = io_inputBit | _GEN_2261; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2263 = _GEN_6085 == 10'h28d ? _GEN_2262 : _GEN_2261; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2264 = ~io_inputBit ? 1'h0 : _GEN_2263; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2265 = _GEN_6085 == 10'h28e ? _GEN_2264 : _GEN_2263; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2266 = io_inputBit | _GEN_2265; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2267 = _GEN_6085 == 10'h28e ? _GEN_2266 : _GEN_2265; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2268 = ~io_inputBit ? 1'h0 : _GEN_2267; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2269 = _GEN_6085 == 10'h28f ? _GEN_2268 : _GEN_2267; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2270 = io_inputBit | _GEN_2269; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2271 = _GEN_6085 == 10'h28f ? _GEN_2270 : _GEN_2269; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2272 = ~io_inputBit ? 1'h0 : _GEN_2271; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2273 = _GEN_6085 == 10'h290 ? _GEN_2272 : _GEN_2271; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2274 = io_inputBit | _GEN_2273; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2275 = _GEN_6085 == 10'h290 ? _GEN_2274 : _GEN_2273; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2276 = ~io_inputBit ? 1'h0 : _GEN_2275; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2277 = _GEN_6085 == 10'h291 ? _GEN_2276 : _GEN_2275; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2278 = io_inputBit | _GEN_2277; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2279 = _GEN_6085 == 10'h291 ? _GEN_2278 : _GEN_2277; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2280 = ~io_inputBit ? 1'h0 : _GEN_2279; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2281 = _GEN_6085 == 10'h292 ? _GEN_2280 : _GEN_2279; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2282 = io_inputBit | _GEN_2281; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2283 = _GEN_6085 == 10'h292 ? _GEN_2282 : _GEN_2281; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2284 = ~io_inputBit ? 1'h0 : _GEN_2283; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2285 = _GEN_6085 == 10'h293 ? _GEN_2284 : _GEN_2283; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2286 = io_inputBit | _GEN_2285; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2287 = _GEN_6085 == 10'h293 ? _GEN_2286 : _GEN_2285; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2288 = ~io_inputBit ? 1'h0 : _GEN_2287; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2289 = _GEN_6085 == 10'h294 ? _GEN_2288 : _GEN_2287; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2290 = io_inputBit | _GEN_2289; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2291 = _GEN_6085 == 10'h294 ? _GEN_2290 : _GEN_2289; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2292 = io_inputBit ? 1'h0 : _GEN_885; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2293 = i == 8'h0 ? _GEN_2292 : _GEN_885; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2294 = ~io_inputBit ? 1'h0 : _GEN_2293; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2295 = i == 8'h1 ? _GEN_2294 : _GEN_2293; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2296 = io_inputBit ? 1'h0 : _GEN_2295; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2297 = i == 8'h4 ? _GEN_2296 : _GEN_2295; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2298 = io_inputBit ? 1'h0 : _GEN_2297; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2299 = i == 8'h9 ? _GEN_2298 : _GEN_2297; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2300 = io_inputBit | _GEN_2299; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2301 = i == 8'h27 ? _GEN_2300 : _GEN_2299; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2302 = io_inputBit ? 1'h0 : _GEN_2301; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2303 = i == 8'h28 ? _GEN_2302 : _GEN_2301; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2304 = ~io_inputBit ? 1'h0 : _GEN_2303; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2305 = i == 8'h4f ? _GEN_2304 : _GEN_2303; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2306 = io_inputBit | _GEN_2305; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2307 = i == 8'h4f ? _GEN_2306 : _GEN_2305; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2308 = ~io_inputBit | _GEN_2307; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2309 = i == 8'h51 ? _GEN_2308 : _GEN_2307; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2310 = ~io_inputBit | _GEN_2309; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2311 = i == 8'ha4 ? _GEN_2310 : _GEN_2309; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2312 = io_inputBit ? 1'h0 : _GEN_2311; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2313 = _GEN_6084 == 9'h14a ? _GEN_2312 : _GEN_2311; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2314 = ~io_inputBit | _GEN_2313; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2315 = _GEN_6085 == 10'h295 ? _GEN_2314 : _GEN_2313; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2316 = io_inputBit ? 1'h0 : _GEN_2315; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2317 = _GEN_6085 == 10'h295 ? _GEN_2316 : _GEN_2315; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2318 = io_inputBit ? 1'h0 : _GEN_963; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2319 = i == 8'h0 ? _GEN_2318 : _GEN_963; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2320 = ~io_inputBit ? 1'h0 : _GEN_2319; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2321 = i == 8'h3 ? _GEN_2320 : _GEN_2319; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2322 = io_inputBit ? 1'h0 : _GEN_2321; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2323 = i == 8'h4 ? _GEN_2322 : _GEN_2321; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2324 = ~io_inputBit ? 1'h0 : _GEN_2323; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2325 = i == 8'h8 ? _GEN_2324 : _GEN_2323; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2326 = io_inputBit ? 1'h0 : _GEN_2325; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2327 = i == 8'h9 ? _GEN_2326 : _GEN_2325; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2328 = ~io_inputBit ? 1'h0 : _GEN_2327; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2329 = i == 8'h12 ? _GEN_2328 : _GEN_2327; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2330 = io_inputBit | _GEN_2329; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2331 = i == 8'h26 ? _GEN_2330 : _GEN_2329; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2332 = io_inputBit ? 1'h0 : _GEN_2331; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2333 = i == 8'h27 ? _GEN_2332 : _GEN_2331; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2334 = io_inputBit ? 1'h0 : _GEN_2333; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2335 = i == 8'h28 ? _GEN_2334 : _GEN_2333; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2336 = ~io_inputBit ? 1'h0 : _GEN_2335; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2337 = i == 8'h4d ? _GEN_2336 : _GEN_2335; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2338 = io_inputBit | _GEN_2337; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2339 = i == 8'h4d ? _GEN_2338 : _GEN_2337; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2340 = ~io_inputBit | _GEN_2339; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2341 = i == 8'h4f ? _GEN_2340 : _GEN_2339; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2342 = io_inputBit ? 1'h0 : _GEN_2341; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2343 = i == 8'h4f ? _GEN_2342 : _GEN_2341; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2344 = ~io_inputBit ? 1'h0 : _GEN_2343; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2345 = i == 8'h51 ? _GEN_2344 : _GEN_2343; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2346 = ~io_inputBit | _GEN_2345; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2347 = i == 8'ha4 ? _GEN_2346 : _GEN_2345; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2348 = io_inputBit ? 1'h0 : _GEN_2347; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2349 = _GEN_6084 == 9'h14a ? _GEN_2348 : _GEN_2347; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2350 = ~io_inputBit | _GEN_2349; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2351 = _GEN_6085 == 10'h295 ? _GEN_2350 : _GEN_2349; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2352 = io_inputBit ? 1'h0 : _GEN_2351; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2353 = _GEN_6085 == 10'h295 ? _GEN_2352 : _GEN_2351; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2354 = io_inputBit ? 1'h0 : _GEN_1083; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2355 = i == 8'h0 ? _GEN_2354 : _GEN_1083; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2356 = ~io_inputBit ? 1'h0 : _GEN_2355; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2357 = i == 8'h3 ? _GEN_2356 : _GEN_2355; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2358 = io_inputBit ? 1'h0 : _GEN_2357; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2359 = i == 8'h4 ? _GEN_2358 : _GEN_2357; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2360 = ~io_inputBit ? 1'h0 : _GEN_2359; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2361 = i == 8'h8 ? _GEN_2360 : _GEN_2359; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2362 = io_inputBit ? 1'h0 : _GEN_2361; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2363 = i == 8'h9 ? _GEN_2362 : _GEN_2361; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2364 = ~io_inputBit ? 1'h0 : _GEN_2363; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2365 = i == 8'h25 ? _GEN_2364 : _GEN_2363; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2366 = io_inputBit ? 1'h0 : _GEN_2365; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2367 = i == 8'h28 ? _GEN_2366 : _GEN_2365; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2368 = ~io_inputBit ? 1'h0 : _GEN_2367; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2369 = i == 8'h4c ? _GEN_2368 : _GEN_2367; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2370 = io_inputBit | _GEN_2369; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2371 = i == 8'h4c ? _GEN_2370 : _GEN_2369; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2372 = ~io_inputBit | _GEN_2371; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2373 = i == 8'h4d ? _GEN_2372 : _GEN_2371; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2374 = io_inputBit ? 1'h0 : _GEN_2373; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2375 = i == 8'h4d ? _GEN_2374 : _GEN_2373; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2376 = ~io_inputBit ? 1'h0 : _GEN_2375; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2377 = i == 8'h4e ? _GEN_2376 : _GEN_2375; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2378 = io_inputBit | _GEN_2377; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2379 = i == 8'h4e ? _GEN_2378 : _GEN_2377; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2380 = ~io_inputBit | _GEN_2379; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2381 = i == 8'h4f ? _GEN_2380 : _GEN_2379; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2382 = io_inputBit ? 1'h0 : _GEN_2381; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2383 = i == 8'h4f ? _GEN_2382 : _GEN_2381; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2384 = ~io_inputBit ? 1'h0 : _GEN_2383; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2385 = i == 8'h50 ? _GEN_2384 : _GEN_2383; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2386 = io_inputBit | _GEN_2385; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2387 = i == 8'h50 ? _GEN_2386 : _GEN_2385; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2388 = ~io_inputBit | _GEN_2387; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2389 = i == 8'h51 ? _GEN_2388 : _GEN_2387; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2390 = io_inputBit ? 1'h0 : _GEN_2389; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2391 = i == 8'h51 ? _GEN_2390 : _GEN_2389; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2392 = io_inputBit ? 1'h0 : _GEN_1273; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2393 = i == 8'h0 ? _GEN_2392 : _GEN_1273; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2394 = ~io_inputBit ? 1'h0 : _GEN_2393; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2395 = i == 8'h3 ? _GEN_2394 : _GEN_2393; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2396 = io_inputBit ? 1'h0 : _GEN_2395; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2397 = i == 8'h4 ? _GEN_2396 : _GEN_2395; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2398 = ~io_inputBit ? 1'h0 : _GEN_2397; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2399 = i == 8'h8 ? _GEN_2398 : _GEN_2397; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2400 = io_inputBit ? 1'h0 : _GEN_2399; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2401 = i == 8'h9 ? _GEN_2400 : _GEN_2399; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2402 = ~io_inputBit ? 1'h0 : _GEN_2401; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2403 = i == 8'h25 ? _GEN_2402 : _GEN_2401; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2404 = io_inputBit ? 1'h0 : _GEN_2403; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2405 = i == 8'h28 ? _GEN_2404 : _GEN_2403; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2406 = ~io_inputBit | _GEN_2405; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2407 = i == 8'h4c ? _GEN_2406 : _GEN_2405; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2408 = io_inputBit ? 1'h0 : _GEN_2407; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2409 = i == 8'h4c ? _GEN_2408 : _GEN_2407; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2410 = ~io_inputBit | _GEN_2409; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2411 = i == 8'h4d ? _GEN_2410 : _GEN_2409; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2412 = io_inputBit ? 1'h0 : _GEN_2411; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2413 = i == 8'h4d ? _GEN_2412 : _GEN_2411; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2414 = ~io_inputBit | _GEN_2413; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2415 = i == 8'h4e ? _GEN_2414 : _GEN_2413; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2416 = io_inputBit ? 1'h0 : _GEN_2415; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2417 = i == 8'h4e ? _GEN_2416 : _GEN_2415; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2418 = ~io_inputBit | _GEN_2417; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2419 = i == 8'h4f ? _GEN_2418 : _GEN_2417; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2420 = io_inputBit ? 1'h0 : _GEN_2419; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2421 = i == 8'h4f ? _GEN_2420 : _GEN_2419; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2422 = ~io_inputBit | _GEN_2421; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2423 = i == 8'h50 ? _GEN_2422 : _GEN_2421; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2424 = io_inputBit ? 1'h0 : _GEN_2423; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2425 = i == 8'h50 ? _GEN_2424 : _GEN_2423; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2426 = ~io_inputBit | _GEN_2425; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2427 = i == 8'h51 ? _GEN_2426 : _GEN_2425; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2428 = io_inputBit ? 1'h0 : _GEN_2427; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2429 = i == 8'h51 ? _GEN_2428 : _GEN_2427; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2430 = io_inputBit ? 1'h0 : _GEN_1545; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2431 = i == 8'h0 ? _GEN_2430 : _GEN_1545; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2432 = ~io_inputBit ? 1'h0 : _GEN_2431; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2433 = i == 8'h3 ? _GEN_2432 : _GEN_2431; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2434 = io_inputBit ? 1'h0 : _GEN_2433; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2435 = i == 8'h4 ? _GEN_2434 : _GEN_2433; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2436 = ~io_inputBit ? 1'h0 : _GEN_2435; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2437 = i == 8'h8 ? _GEN_2436 : _GEN_2435; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2438 = io_inputBit ? 1'h0 : _GEN_2437; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2439 = i == 8'h9 ? _GEN_2438 : _GEN_2437; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2440 = io_inputBit ? 1'h0 : _GEN_2439; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2441 = i == 8'h28 ? _GEN_2440 : _GEN_2439; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2442 = ~io_inputBit ? 1'h0 : _GEN_2441; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2443 = i == 8'h4b ? _GEN_2442 : _GEN_2441; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2444 = ~io_inputBit ? 1'h0 : _GEN_2443; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2445 = i == 8'h98 ? _GEN_2444 : _GEN_2443; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2446 = io_inputBit | _GEN_2445; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2447 = i == 8'h98 ? _GEN_2446 : _GEN_2445; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2448 = ~io_inputBit ? 1'h0 : _GEN_2447; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2449 = i == 8'h99 ? _GEN_2448 : _GEN_2447; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2450 = io_inputBit | _GEN_2449; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2451 = i == 8'h99 ? _GEN_2450 : _GEN_2449; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2452 = ~io_inputBit ? 1'h0 : _GEN_2451; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2453 = i == 8'h9a ? _GEN_2452 : _GEN_2451; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2454 = io_inputBit | _GEN_2453; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2455 = i == 8'h9a ? _GEN_2454 : _GEN_2453; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2456 = ~io_inputBit ? 1'h0 : _GEN_2455; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2457 = i == 8'h9b ? _GEN_2456 : _GEN_2455; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2458 = io_inputBit | _GEN_2457; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2459 = i == 8'h9b ? _GEN_2458 : _GEN_2457; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2460 = ~io_inputBit ? 1'h0 : _GEN_2459; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2461 = i == 8'h9c ? _GEN_2460 : _GEN_2459; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2462 = io_inputBit | _GEN_2461; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2463 = i == 8'h9c ? _GEN_2462 : _GEN_2461; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2464 = ~io_inputBit ? 1'h0 : _GEN_2463; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2465 = i == 8'h9d ? _GEN_2464 : _GEN_2463; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2466 = io_inputBit | _GEN_2465; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2467 = i == 8'h9d ? _GEN_2466 : _GEN_2465; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2468 = ~io_inputBit ? 1'h0 : _GEN_2467; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2469 = i == 8'h9e ? _GEN_2468 : _GEN_2467; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2470 = io_inputBit | _GEN_2469; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2471 = i == 8'h9e ? _GEN_2470 : _GEN_2469; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2472 = ~io_inputBit ? 1'h0 : _GEN_2471; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2473 = i == 8'h9f ? _GEN_2472 : _GEN_2471; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2474 = io_inputBit | _GEN_2473; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2475 = i == 8'h9f ? _GEN_2474 : _GEN_2473; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2476 = ~io_inputBit ? 1'h0 : _GEN_2475; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2477 = i == 8'ha0 ? _GEN_2476 : _GEN_2475; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2478 = io_inputBit | _GEN_2477; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2479 = i == 8'ha0 ? _GEN_2478 : _GEN_2477; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2480 = ~io_inputBit ? 1'h0 : _GEN_2479; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2481 = i == 8'ha1 ? _GEN_2480 : _GEN_2479; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2482 = io_inputBit | _GEN_2481; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2483 = i == 8'ha1 ? _GEN_2482 : _GEN_2481; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2484 = ~io_inputBit ? 1'h0 : _GEN_2483; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2485 = i == 8'ha2 ? _GEN_2484 : _GEN_2483; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2486 = io_inputBit | _GEN_2485; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2487 = i == 8'ha2 ? _GEN_2486 : _GEN_2485; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2488 = ~io_inputBit ? 1'h0 : _GEN_2487; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2489 = i == 8'ha3 ? _GEN_2488 : _GEN_2487; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2490 = io_inputBit | _GEN_2489; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2491 = i == 8'ha3 ? _GEN_2490 : _GEN_2489; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2492 = ~io_inputBit ? 1'h0 : _GEN_2491; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2493 = i == 8'ha4 ? _GEN_2492 : _GEN_2491; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2494 = io_inputBit ? 1'h0 : _GEN_2493; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2495 = _GEN_6084 == 9'h14a ? _GEN_2494 : _GEN_2493; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2496 = ~io_inputBit | _GEN_2495; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2497 = _GEN_6085 == 10'h295 ? _GEN_2496 : _GEN_2495; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2498 = io_inputBit ? 1'h0 : _GEN_2497; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2499 = _GEN_6085 == 10'h295 ? _GEN_2498 : _GEN_2497; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2500 = io_inputBit ? 1'h0 : _GEN_1867; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2501 = i == 8'h0 ? _GEN_2500 : _GEN_1867; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2502 = ~io_inputBit ? 1'h0 : _GEN_2501; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2503 = i == 8'h3 ? _GEN_2502 : _GEN_2501; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2504 = io_inputBit ? 1'h0 : _GEN_2503; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2505 = i == 8'h4 ? _GEN_2504 : _GEN_2503; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2506 = ~io_inputBit ? 1'h0 : _GEN_2505; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2507 = i == 8'h8 ? _GEN_2506 : _GEN_2505; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2508 = io_inputBit ? 1'h0 : _GEN_2507; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2509 = i == 8'h9 ? _GEN_2508 : _GEN_2507; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2510 = io_inputBit ? 1'h0 : _GEN_2509; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2511 = i == 8'h28 ? _GEN_2510 : _GEN_2509; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2512 = ~io_inputBit ? 1'h0 : _GEN_2511; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2513 = i == 8'h4b ? _GEN_2512 : _GEN_2511; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2514 = io_inputBit ? 1'h0 : _GEN_2513; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2515 = i == 8'ha4 ? _GEN_2514 : _GEN_2513; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2516 = ~io_inputBit ? 1'h0 : _GEN_2515; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2517 = _GEN_6084 == 9'h131 ? _GEN_2516 : _GEN_2515; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2518 = io_inputBit | _GEN_2517; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2519 = _GEN_6084 == 9'h131 ? _GEN_2518 : _GEN_2517; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2520 = ~io_inputBit ? 1'h0 : _GEN_2519; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2521 = _GEN_6084 == 9'h132 ? _GEN_2520 : _GEN_2519; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2522 = io_inputBit | _GEN_2521; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2523 = _GEN_6084 == 9'h132 ? _GEN_2522 : _GEN_2521; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2524 = ~io_inputBit ? 1'h0 : _GEN_2523; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2525 = _GEN_6084 == 9'h133 ? _GEN_2524 : _GEN_2523; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2526 = io_inputBit | _GEN_2525; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2527 = _GEN_6084 == 9'h133 ? _GEN_2526 : _GEN_2525; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2528 = ~io_inputBit ? 1'h0 : _GEN_2527; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2529 = _GEN_6084 == 9'h134 ? _GEN_2528 : _GEN_2527; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2530 = io_inputBit | _GEN_2529; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2531 = _GEN_6084 == 9'h134 ? _GEN_2530 : _GEN_2529; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2532 = ~io_inputBit ? 1'h0 : _GEN_2531; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2533 = _GEN_6084 == 9'h135 ? _GEN_2532 : _GEN_2531; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2534 = io_inputBit | _GEN_2533; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2535 = _GEN_6084 == 9'h135 ? _GEN_2534 : _GEN_2533; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2536 = ~io_inputBit ? 1'h0 : _GEN_2535; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2537 = _GEN_6084 == 9'h136 ? _GEN_2536 : _GEN_2535; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2538 = io_inputBit | _GEN_2537; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2539 = _GEN_6084 == 9'h136 ? _GEN_2538 : _GEN_2537; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2540 = ~io_inputBit ? 1'h0 : _GEN_2539; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2541 = _GEN_6084 == 9'h137 ? _GEN_2540 : _GEN_2539; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2542 = io_inputBit | _GEN_2541; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2543 = _GEN_6084 == 9'h137 ? _GEN_2542 : _GEN_2541; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2544 = ~io_inputBit ? 1'h0 : _GEN_2543; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2545 = _GEN_6084 == 9'h138 ? _GEN_2544 : _GEN_2543; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2546 = io_inputBit | _GEN_2545; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2547 = _GEN_6084 == 9'h138 ? _GEN_2546 : _GEN_2545; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2548 = ~io_inputBit ? 1'h0 : _GEN_2547; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2549 = _GEN_6084 == 9'h139 ? _GEN_2548 : _GEN_2547; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2550 = io_inputBit | _GEN_2549; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2551 = _GEN_6084 == 9'h139 ? _GEN_2550 : _GEN_2549; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2552 = ~io_inputBit ? 1'h0 : _GEN_2551; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2553 = _GEN_6084 == 9'h13a ? _GEN_2552 : _GEN_2551; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2554 = io_inputBit | _GEN_2553; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2555 = _GEN_6084 == 9'h13a ? _GEN_2554 : _GEN_2553; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2556 = ~io_inputBit ? 1'h0 : _GEN_2555; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2557 = _GEN_6084 == 9'h13b ? _GEN_2556 : _GEN_2555; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2558 = io_inputBit | _GEN_2557; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2559 = _GEN_6084 == 9'h13b ? _GEN_2558 : _GEN_2557; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2560 = ~io_inputBit ? 1'h0 : _GEN_2559; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2561 = _GEN_6084 == 9'h13c ? _GEN_2560 : _GEN_2559; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2562 = io_inputBit | _GEN_2561; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2563 = _GEN_6084 == 9'h13c ? _GEN_2562 : _GEN_2561; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2564 = ~io_inputBit ? 1'h0 : _GEN_2563; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2565 = _GEN_6084 == 9'h13d ? _GEN_2564 : _GEN_2563; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2566 = io_inputBit | _GEN_2565; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2567 = _GEN_6084 == 9'h13d ? _GEN_2566 : _GEN_2565; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2568 = ~io_inputBit ? 1'h0 : _GEN_2567; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2569 = _GEN_6084 == 9'h13e ? _GEN_2568 : _GEN_2567; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2570 = io_inputBit | _GEN_2569; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2571 = _GEN_6084 == 9'h13e ? _GEN_2570 : _GEN_2569; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2572 = ~io_inputBit ? 1'h0 : _GEN_2571; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2573 = _GEN_6084 == 9'h13f ? _GEN_2572 : _GEN_2571; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2574 = io_inputBit | _GEN_2573; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2575 = _GEN_6084 == 9'h13f ? _GEN_2574 : _GEN_2573; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2576 = ~io_inputBit ? 1'h0 : _GEN_2575; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2577 = _GEN_6084 == 9'h140 ? _GEN_2576 : _GEN_2575; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2578 = io_inputBit | _GEN_2577; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2579 = _GEN_6084 == 9'h140 ? _GEN_2578 : _GEN_2577; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2580 = ~io_inputBit ? 1'h0 : _GEN_2579; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2581 = _GEN_6084 == 9'h141 ? _GEN_2580 : _GEN_2579; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2582 = io_inputBit | _GEN_2581; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2583 = _GEN_6084 == 9'h141 ? _GEN_2582 : _GEN_2581; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2584 = ~io_inputBit ? 1'h0 : _GEN_2583; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2585 = _GEN_6084 == 9'h142 ? _GEN_2584 : _GEN_2583; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2586 = io_inputBit | _GEN_2585; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2587 = _GEN_6084 == 9'h142 ? _GEN_2586 : _GEN_2585; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2588 = ~io_inputBit ? 1'h0 : _GEN_2587; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2589 = _GEN_6084 == 9'h143 ? _GEN_2588 : _GEN_2587; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2590 = io_inputBit | _GEN_2589; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2591 = _GEN_6084 == 9'h143 ? _GEN_2590 : _GEN_2589; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2592 = ~io_inputBit ? 1'h0 : _GEN_2591; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2593 = _GEN_6084 == 9'h144 ? _GEN_2592 : _GEN_2591; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2594 = io_inputBit | _GEN_2593; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2595 = _GEN_6084 == 9'h144 ? _GEN_2594 : _GEN_2593; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2596 = ~io_inputBit ? 1'h0 : _GEN_2595; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2597 = _GEN_6084 == 9'h145 ? _GEN_2596 : _GEN_2595; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2598 = io_inputBit | _GEN_2597; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2599 = _GEN_6084 == 9'h145 ? _GEN_2598 : _GEN_2597; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2600 = ~io_inputBit ? 1'h0 : _GEN_2599; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2601 = _GEN_6084 == 9'h146 ? _GEN_2600 : _GEN_2599; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2602 = io_inputBit | _GEN_2601; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2603 = _GEN_6084 == 9'h146 ? _GEN_2602 : _GEN_2601; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2604 = ~io_inputBit ? 1'h0 : _GEN_2603; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2605 = _GEN_6084 == 9'h147 ? _GEN_2604 : _GEN_2603; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2606 = io_inputBit | _GEN_2605; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2607 = _GEN_6084 == 9'h147 ? _GEN_2606 : _GEN_2605; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2608 = ~io_inputBit ? 1'h0 : _GEN_2607; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2609 = _GEN_6084 == 9'h148 ? _GEN_2608 : _GEN_2607; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2610 = io_inputBit | _GEN_2609; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2611 = _GEN_6084 == 9'h148 ? _GEN_2610 : _GEN_2609; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2612 = ~io_inputBit ? 1'h0 : _GEN_2611; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2613 = _GEN_6084 == 9'h149 ? _GEN_2612 : _GEN_2611; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2614 = io_inputBit | _GEN_2613; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2615 = _GEN_6084 == 9'h149 ? _GEN_2614 : _GEN_2613; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2616 = io_inputBit ? 1'h0 : _GEN_2291; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2617 = i == 8'h0 ? _GEN_2616 : _GEN_2291; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2618 = ~io_inputBit ? 1'h0 : _GEN_2617; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2619 = i == 8'h3 ? _GEN_2618 : _GEN_2617; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2620 = io_inputBit ? 1'h0 : _GEN_2619; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2621 = i == 8'h4 ? _GEN_2620 : _GEN_2619; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2622 = ~io_inputBit ? 1'h0 : _GEN_2621; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2623 = i == 8'h8 ? _GEN_2622 : _GEN_2621; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2624 = io_inputBit ? 1'h0 : _GEN_2623; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2625 = i == 8'h9 ? _GEN_2624 : _GEN_2623; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2626 = io_inputBit ? 1'h0 : _GEN_2625; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2627 = i == 8'h28 ? _GEN_2626 : _GEN_2625; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2628 = ~io_inputBit ? 1'h0 : _GEN_2627; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2629 = i == 8'h4b ? _GEN_2628 : _GEN_2627; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2630 = io_inputBit ? 1'h0 : _GEN_2629; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2631 = i == 8'ha4 ? _GEN_2630 : _GEN_2629; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2632 = ~io_inputBit ? 1'h0 : _GEN_2631; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2633 = _GEN_6085 == 10'h263 ? _GEN_2632 : _GEN_2631; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2634 = io_inputBit | _GEN_2633; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2635 = _GEN_6085 == 10'h263 ? _GEN_2634 : _GEN_2633; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2636 = ~io_inputBit ? 1'h0 : _GEN_2635; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2637 = _GEN_6085 == 10'h264 ? _GEN_2636 : _GEN_2635; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2638 = io_inputBit | _GEN_2637; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2639 = _GEN_6085 == 10'h264 ? _GEN_2638 : _GEN_2637; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2640 = ~io_inputBit ? 1'h0 : _GEN_2639; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2641 = _GEN_6085 == 10'h265 ? _GEN_2640 : _GEN_2639; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2642 = io_inputBit | _GEN_2641; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2643 = _GEN_6085 == 10'h265 ? _GEN_2642 : _GEN_2641; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2644 = ~io_inputBit ? 1'h0 : _GEN_2643; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2645 = _GEN_6085 == 10'h266 ? _GEN_2644 : _GEN_2643; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2646 = io_inputBit | _GEN_2645; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2647 = _GEN_6085 == 10'h266 ? _GEN_2646 : _GEN_2645; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2648 = ~io_inputBit ? 1'h0 : _GEN_2647; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2649 = _GEN_6085 == 10'h267 ? _GEN_2648 : _GEN_2647; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2650 = io_inputBit | _GEN_2649; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2651 = _GEN_6085 == 10'h267 ? _GEN_2650 : _GEN_2649; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2652 = ~io_inputBit ? 1'h0 : _GEN_2651; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2653 = _GEN_6085 == 10'h268 ? _GEN_2652 : _GEN_2651; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2654 = io_inputBit | _GEN_2653; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2655 = _GEN_6085 == 10'h268 ? _GEN_2654 : _GEN_2653; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2656 = ~io_inputBit ? 1'h0 : _GEN_2655; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2657 = _GEN_6085 == 10'h269 ? _GEN_2656 : _GEN_2655; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2658 = io_inputBit | _GEN_2657; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2659 = _GEN_6085 == 10'h269 ? _GEN_2658 : _GEN_2657; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2660 = ~io_inputBit ? 1'h0 : _GEN_2659; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2661 = _GEN_6085 == 10'h26a ? _GEN_2660 : _GEN_2659; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2662 = io_inputBit | _GEN_2661; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2663 = _GEN_6085 == 10'h26a ? _GEN_2662 : _GEN_2661; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2664 = ~io_inputBit ? 1'h0 : _GEN_2663; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2665 = _GEN_6085 == 10'h26b ? _GEN_2664 : _GEN_2663; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2666 = io_inputBit | _GEN_2665; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2667 = _GEN_6085 == 10'h26b ? _GEN_2666 : _GEN_2665; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2668 = ~io_inputBit ? 1'h0 : _GEN_2667; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2669 = _GEN_6085 == 10'h26c ? _GEN_2668 : _GEN_2667; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2670 = io_inputBit | _GEN_2669; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2671 = _GEN_6085 == 10'h26c ? _GEN_2670 : _GEN_2669; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2672 = ~io_inputBit ? 1'h0 : _GEN_2671; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2673 = _GEN_6085 == 10'h26d ? _GEN_2672 : _GEN_2671; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2674 = io_inputBit | _GEN_2673; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2675 = _GEN_6085 == 10'h26d ? _GEN_2674 : _GEN_2673; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2676 = ~io_inputBit ? 1'h0 : _GEN_2675; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2677 = _GEN_6085 == 10'h26e ? _GEN_2676 : _GEN_2675; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2678 = io_inputBit | _GEN_2677; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2679 = _GEN_6085 == 10'h26e ? _GEN_2678 : _GEN_2677; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2680 = ~io_inputBit ? 1'h0 : _GEN_2679; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2681 = _GEN_6085 == 10'h26f ? _GEN_2680 : _GEN_2679; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2682 = io_inputBit | _GEN_2681; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2683 = _GEN_6085 == 10'h26f ? _GEN_2682 : _GEN_2681; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2684 = ~io_inputBit ? 1'h0 : _GEN_2683; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2685 = _GEN_6085 == 10'h270 ? _GEN_2684 : _GEN_2683; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2686 = io_inputBit | _GEN_2685; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2687 = _GEN_6085 == 10'h270 ? _GEN_2686 : _GEN_2685; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2688 = ~io_inputBit ? 1'h0 : _GEN_2687; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2689 = _GEN_6085 == 10'h271 ? _GEN_2688 : _GEN_2687; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2690 = io_inputBit | _GEN_2689; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2691 = _GEN_6085 == 10'h271 ? _GEN_2690 : _GEN_2689; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2692 = ~io_inputBit ? 1'h0 : _GEN_2691; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2693 = _GEN_6085 == 10'h272 ? _GEN_2692 : _GEN_2691; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2694 = io_inputBit | _GEN_2693; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2695 = _GEN_6085 == 10'h272 ? _GEN_2694 : _GEN_2693; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2696 = ~io_inputBit ? 1'h0 : _GEN_2695; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2697 = _GEN_6085 == 10'h273 ? _GEN_2696 : _GEN_2695; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2698 = io_inputBit | _GEN_2697; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2699 = _GEN_6085 == 10'h273 ? _GEN_2698 : _GEN_2697; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2700 = ~io_inputBit ? 1'h0 : _GEN_2699; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2701 = _GEN_6085 == 10'h274 ? _GEN_2700 : _GEN_2699; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2702 = io_inputBit | _GEN_2701; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2703 = _GEN_6085 == 10'h274 ? _GEN_2702 : _GEN_2701; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2704 = ~io_inputBit ? 1'h0 : _GEN_2703; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2705 = _GEN_6085 == 10'h275 ? _GEN_2704 : _GEN_2703; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2706 = io_inputBit | _GEN_2705; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2707 = _GEN_6085 == 10'h275 ? _GEN_2706 : _GEN_2705; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2708 = ~io_inputBit ? 1'h0 : _GEN_2707; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2709 = _GEN_6085 == 10'h276 ? _GEN_2708 : _GEN_2707; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2710 = io_inputBit | _GEN_2709; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2711 = _GEN_6085 == 10'h276 ? _GEN_2710 : _GEN_2709; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2712 = ~io_inputBit ? 1'h0 : _GEN_2711; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2713 = _GEN_6085 == 10'h277 ? _GEN_2712 : _GEN_2711; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2714 = io_inputBit | _GEN_2713; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2715 = _GEN_6085 == 10'h277 ? _GEN_2714 : _GEN_2713; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2716 = ~io_inputBit ? 1'h0 : _GEN_2715; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2717 = _GEN_6085 == 10'h278 ? _GEN_2716 : _GEN_2715; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2718 = io_inputBit | _GEN_2717; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2719 = _GEN_6085 == 10'h278 ? _GEN_2718 : _GEN_2717; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2720 = ~io_inputBit ? 1'h0 : _GEN_2719; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2721 = _GEN_6085 == 10'h279 ? _GEN_2720 : _GEN_2719; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2722 = io_inputBit | _GEN_2721; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2723 = _GEN_6085 == 10'h279 ? _GEN_2722 : _GEN_2721; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2724 = ~io_inputBit ? 1'h0 : _GEN_2723; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2725 = _GEN_6085 == 10'h27a ? _GEN_2724 : _GEN_2723; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2726 = io_inputBit | _GEN_2725; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2727 = _GEN_6085 == 10'h27a ? _GEN_2726 : _GEN_2725; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2728 = ~io_inputBit ? 1'h0 : _GEN_2727; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2729 = _GEN_6085 == 10'h27b ? _GEN_2728 : _GEN_2727; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2730 = io_inputBit | _GEN_2729; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2731 = _GEN_6085 == 10'h27b ? _GEN_2730 : _GEN_2729; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2732 = ~io_inputBit ? 1'h0 : _GEN_2731; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2733 = _GEN_6085 == 10'h27c ? _GEN_2732 : _GEN_2731; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2734 = io_inputBit | _GEN_2733; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2735 = _GEN_6085 == 10'h27c ? _GEN_2734 : _GEN_2733; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2736 = ~io_inputBit ? 1'h0 : _GEN_2735; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2737 = _GEN_6085 == 10'h27d ? _GEN_2736 : _GEN_2735; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2738 = io_inputBit | _GEN_2737; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2739 = _GEN_6085 == 10'h27d ? _GEN_2738 : _GEN_2737; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2740 = ~io_inputBit ? 1'h0 : _GEN_2739; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2741 = _GEN_6085 == 10'h27e ? _GEN_2740 : _GEN_2739; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2742 = io_inputBit | _GEN_2741; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2743 = _GEN_6085 == 10'h27e ? _GEN_2742 : _GEN_2741; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2744 = ~io_inputBit ? 1'h0 : _GEN_2743; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2745 = _GEN_6085 == 10'h27f ? _GEN_2744 : _GEN_2743; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2746 = io_inputBit | _GEN_2745; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2747 = _GEN_6085 == 10'h27f ? _GEN_2746 : _GEN_2745; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2748 = ~io_inputBit ? 1'h0 : _GEN_2747; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2749 = _GEN_6085 == 10'h280 ? _GEN_2748 : _GEN_2747; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2750 = io_inputBit | _GEN_2749; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2751 = _GEN_6085 == 10'h280 ? _GEN_2750 : _GEN_2749; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2752 = ~io_inputBit ? 1'h0 : _GEN_2751; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2753 = _GEN_6085 == 10'h281 ? _GEN_2752 : _GEN_2751; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2754 = io_inputBit | _GEN_2753; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2755 = _GEN_6085 == 10'h281 ? _GEN_2754 : _GEN_2753; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2756 = ~io_inputBit ? 1'h0 : _GEN_2755; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2757 = _GEN_6085 == 10'h282 ? _GEN_2756 : _GEN_2755; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2758 = io_inputBit | _GEN_2757; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2759 = _GEN_6085 == 10'h282 ? _GEN_2758 : _GEN_2757; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2760 = ~io_inputBit ? 1'h0 : _GEN_2759; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2761 = _GEN_6085 == 10'h283 ? _GEN_2760 : _GEN_2759; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2762 = io_inputBit | _GEN_2761; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2763 = _GEN_6085 == 10'h283 ? _GEN_2762 : _GEN_2761; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2764 = ~io_inputBit ? 1'h0 : _GEN_2763; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2765 = _GEN_6085 == 10'h284 ? _GEN_2764 : _GEN_2763; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2766 = io_inputBit | _GEN_2765; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2767 = _GEN_6085 == 10'h284 ? _GEN_2766 : _GEN_2765; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2768 = ~io_inputBit ? 1'h0 : _GEN_2767; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2769 = _GEN_6085 == 10'h285 ? _GEN_2768 : _GEN_2767; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2770 = io_inputBit | _GEN_2769; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2771 = _GEN_6085 == 10'h285 ? _GEN_2770 : _GEN_2769; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2772 = ~io_inputBit ? 1'h0 : _GEN_2771; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2773 = _GEN_6085 == 10'h286 ? _GEN_2772 : _GEN_2771; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2774 = io_inputBit | _GEN_2773; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2775 = _GEN_6085 == 10'h286 ? _GEN_2774 : _GEN_2773; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2776 = ~io_inputBit ? 1'h0 : _GEN_2775; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2777 = _GEN_6085 == 10'h287 ? _GEN_2776 : _GEN_2775; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2778 = io_inputBit | _GEN_2777; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2779 = _GEN_6085 == 10'h287 ? _GEN_2778 : _GEN_2777; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2780 = ~io_inputBit ? 1'h0 : _GEN_2779; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2781 = _GEN_6085 == 10'h288 ? _GEN_2780 : _GEN_2779; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2782 = io_inputBit | _GEN_2781; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2783 = _GEN_6085 == 10'h288 ? _GEN_2782 : _GEN_2781; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2784 = ~io_inputBit ? 1'h0 : _GEN_2783; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2785 = _GEN_6085 == 10'h289 ? _GEN_2784 : _GEN_2783; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2786 = io_inputBit | _GEN_2785; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2787 = _GEN_6085 == 10'h289 ? _GEN_2786 : _GEN_2785; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2788 = ~io_inputBit ? 1'h0 : _GEN_2787; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2789 = _GEN_6085 == 10'h28a ? _GEN_2788 : _GEN_2787; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2790 = io_inputBit | _GEN_2789; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2791 = _GEN_6085 == 10'h28a ? _GEN_2790 : _GEN_2789; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2792 = ~io_inputBit ? 1'h0 : _GEN_2791; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2793 = _GEN_6085 == 10'h28b ? _GEN_2792 : _GEN_2791; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2794 = io_inputBit | _GEN_2793; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2795 = _GEN_6085 == 10'h28b ? _GEN_2794 : _GEN_2793; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2796 = ~io_inputBit ? 1'h0 : _GEN_2795; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2797 = _GEN_6085 == 10'h28c ? _GEN_2796 : _GEN_2795; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2798 = io_inputBit | _GEN_2797; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2799 = _GEN_6085 == 10'h28c ? _GEN_2798 : _GEN_2797; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2800 = ~io_inputBit ? 1'h0 : _GEN_2799; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2801 = _GEN_6085 == 10'h28d ? _GEN_2800 : _GEN_2799; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2802 = io_inputBit | _GEN_2801; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2803 = _GEN_6085 == 10'h28d ? _GEN_2802 : _GEN_2801; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2804 = ~io_inputBit ? 1'h0 : _GEN_2803; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2805 = _GEN_6085 == 10'h28e ? _GEN_2804 : _GEN_2803; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2806 = io_inputBit | _GEN_2805; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2807 = _GEN_6085 == 10'h28e ? _GEN_2806 : _GEN_2805; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2808 = ~io_inputBit ? 1'h0 : _GEN_2807; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2809 = _GEN_6085 == 10'h28f ? _GEN_2808 : _GEN_2807; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2810 = io_inputBit | _GEN_2809; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2811 = _GEN_6085 == 10'h28f ? _GEN_2810 : _GEN_2809; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2812 = ~io_inputBit ? 1'h0 : _GEN_2811; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2813 = _GEN_6085 == 10'h290 ? _GEN_2812 : _GEN_2811; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2814 = io_inputBit | _GEN_2813; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2815 = _GEN_6085 == 10'h290 ? _GEN_2814 : _GEN_2813; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2816 = ~io_inputBit ? 1'h0 : _GEN_2815; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2817 = _GEN_6085 == 10'h291 ? _GEN_2816 : _GEN_2815; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2818 = io_inputBit | _GEN_2817; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2819 = _GEN_6085 == 10'h291 ? _GEN_2818 : _GEN_2817; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2820 = ~io_inputBit ? 1'h0 : _GEN_2819; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2821 = _GEN_6085 == 10'h292 ? _GEN_2820 : _GEN_2819; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2822 = io_inputBit | _GEN_2821; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2823 = _GEN_6085 == 10'h292 ? _GEN_2822 : _GEN_2821; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2824 = ~io_inputBit ? 1'h0 : _GEN_2823; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2825 = _GEN_6085 == 10'h293 ? _GEN_2824 : _GEN_2823; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2826 = io_inputBit | _GEN_2825; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2827 = _GEN_6085 == 10'h293 ? _GEN_2826 : _GEN_2825; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2828 = ~io_inputBit ? 1'h0 : _GEN_2827; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2829 = _GEN_6085 == 10'h294 ? _GEN_2828 : _GEN_2827; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2830 = io_inputBit | _GEN_2829; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2831 = _GEN_6085 == 10'h294 ? _GEN_2830 : _GEN_2829; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2832 = io_inputBit ? 1'h0 : _GEN_2317; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2833 = i == 8'h0 ? _GEN_2832 : _GEN_2317; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2834 = ~io_inputBit ? 1'h0 : _GEN_2833; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2835 = i == 8'h1 ? _GEN_2834 : _GEN_2833; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2836 = ~io_inputBit ? 1'h0 : _GEN_2835; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2837 = i == 8'h4 ? _GEN_2836 : _GEN_2835; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2838 = io_inputBit | _GEN_2837; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2839 = i == 8'h15 ? _GEN_2838 : _GEN_2837; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2840 = ~io_inputBit | _GEN_2839; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2841 = i == 8'h16 ? _GEN_2840 : _GEN_2839; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2842 = ~io_inputBit ? 1'h0 : _GEN_2841; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2843 = i == 8'h2b ? _GEN_2842 : _GEN_2841; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2844 = io_inputBit ? 1'h0 : _GEN_2843; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2845 = i == 8'h2e ? _GEN_2844 : _GEN_2843; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2846 = ~io_inputBit ? 1'h0 : _GEN_2845; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2847 = i == 8'h58 ? _GEN_2846 : _GEN_2845; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2848 = io_inputBit ? 1'h0 : _GEN_2847; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2849 = i == 8'h5d ? _GEN_2848 : _GEN_2847; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2850 = ~io_inputBit ? 1'h0 : _GEN_2849; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2851 = i == 8'hb2 ? _GEN_2850 : _GEN_2849; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2852 = ~io_inputBit | _GEN_2851; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2853 = i == 8'hbb ? _GEN_2852 : _GEN_2851; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2854 = ~io_inputBit ? 1'h0 : _GEN_2853; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2855 = _GEN_6084 == 9'h166 ? _GEN_2854 : _GEN_2853; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2856 = io_inputBit | _GEN_2855; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2857 = _GEN_6084 == 9'h166 ? _GEN_2856 : _GEN_2855; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2858 = ~io_inputBit | _GEN_2857; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2859 = _GEN_6084 == 9'h178 ? _GEN_2858 : _GEN_2857; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2860 = ~io_inputBit | _GEN_2859; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2861 = _GEN_6085 == 10'h2f2 ? _GEN_2860 : _GEN_2859; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2862 = io_inputBit ? 1'h0 : _GEN_2861; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2863 = _GEN_6085 == 10'h2f2 ? _GEN_2862 : _GEN_2861; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2864 = ~io_inputBit ? 1'h0 : _GEN_2353; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2865 = i == 8'h1 ? _GEN_2864 : _GEN_2353; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2866 = io_inputBit ? 1'h0 : _GEN_2865; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2867 = i == 8'h2 ? _GEN_2866 : _GEN_2865; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2868 = io_inputBit ? 1'h0 : _GEN_2867; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2869 = i == 8'h5 ? _GEN_2868 : _GEN_2867; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2870 = ~io_inputBit ? 1'h0 : _GEN_2869; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2871 = i == 8'h9 ? _GEN_2870 : _GEN_2869; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2872 = io_inputBit ? 1'h0 : _GEN_2871; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2873 = i == 8'hb ? _GEN_2872 : _GEN_2871; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2874 = ~io_inputBit ? 1'h0 : _GEN_2873; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2875 = i == 8'h14 ? _GEN_2874 : _GEN_2873; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2876 = io_inputBit ? 1'h0 : _GEN_2875; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2877 = i == 8'h17 ? _GEN_2876 : _GEN_2875; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2878 = ~io_inputBit ? 1'h0 : _GEN_2877; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2879 = i == 8'h2a ? _GEN_2878 : _GEN_2877; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2880 = ~io_inputBit | _GEN_2879; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2881 = i == 8'h2b ? _GEN_2880 : _GEN_2879; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2882 = ~io_inputBit ? 1'h0 : _GEN_2881; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2883 = i == 8'h2c ? _GEN_2882 : _GEN_2881; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2884 = io_inputBit ? 1'h0 : _GEN_2883; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2885 = i == 8'h2d ? _GEN_2884 : _GEN_2883; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2886 = io_inputBit | _GEN_2885; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2887 = i == 8'h2e ? _GEN_2886 : _GEN_2885; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2888 = io_inputBit ? 1'h0 : _GEN_2887; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2889 = i == 8'h2f ? _GEN_2888 : _GEN_2887; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2890 = ~io_inputBit ? 1'h0 : _GEN_2889; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2891 = i == 8'h56 ? _GEN_2890 : _GEN_2889; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2892 = ~io_inputBit | _GEN_2891; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2893 = i == 8'h58 ? _GEN_2892 : _GEN_2891; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2894 = ~io_inputBit ? 1'h0 : _GEN_2893; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2895 = i == 8'h5a ? _GEN_2894 : _GEN_2893; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2896 = io_inputBit ? 1'h0 : _GEN_2895; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2897 = i == 8'h5b ? _GEN_2896 : _GEN_2895; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2898 = io_inputBit | _GEN_2897; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2899 = i == 8'h5d ? _GEN_2898 : _GEN_2897; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2900 = io_inputBit ? 1'h0 : _GEN_2899; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2901 = i == 8'h5f ? _GEN_2900 : _GEN_2899; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2902 = ~io_inputBit ? 1'h0 : _GEN_2901; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2903 = i == 8'hae ? _GEN_2902 : _GEN_2901; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2904 = ~io_inputBit | _GEN_2903; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2905 = i == 8'hb2 ? _GEN_2904 : _GEN_2903; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2906 = ~io_inputBit ? 1'h0 : _GEN_2905; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2907 = i == 8'hb6 ? _GEN_2906 : _GEN_2905; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2908 = ~io_inputBit | _GEN_2907; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2909 = i == 8'hb7 ? _GEN_2908 : _GEN_2907; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2910 = ~io_inputBit ? 1'h0 : _GEN_2909; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2911 = i == 8'hbb ? _GEN_2910 : _GEN_2909; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2912 = ~io_inputBit | _GEN_2911; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2913 = i == 8'hbf ? _GEN_2912 : _GEN_2911; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2914 = ~io_inputBit ? 1'h0 : _GEN_2913; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2915 = _GEN_6084 == 9'h15e ? _GEN_2914 : _GEN_2913; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2916 = io_inputBit | _GEN_2915; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2917 = _GEN_6084 == 9'h15e ? _GEN_2916 : _GEN_2915; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2918 = ~io_inputBit | _GEN_2917; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2919 = _GEN_6084 == 9'h166 ? _GEN_2918 : _GEN_2917; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2920 = io_inputBit ? 1'h0 : _GEN_2919; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2921 = _GEN_6084 == 9'h166 ? _GEN_2920 : _GEN_2919; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2922 = ~io_inputBit ? 1'h0 : _GEN_2921; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2923 = _GEN_6084 == 9'h16e ? _GEN_2922 : _GEN_2921; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2924 = io_inputBit | _GEN_2923; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2925 = _GEN_6084 == 9'h16e ? _GEN_2924 : _GEN_2923; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2926 = ~io_inputBit | _GEN_2925; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2927 = _GEN_6084 == 9'h170 ? _GEN_2926 : _GEN_2925; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2928 = ~io_inputBit ? 1'h0 : _GEN_2927; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2929 = _GEN_6084 == 9'h178 ? _GEN_2928 : _GEN_2927; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2930 = ~io_inputBit | _GEN_2929; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2931 = _GEN_6084 == 9'h180 ? _GEN_2930 : _GEN_2929; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2932 = ~io_inputBit | _GEN_2931; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2933 = _GEN_6085 == 10'h2e2 ? _GEN_2932 : _GEN_2931; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2934 = io_inputBit ? 1'h0 : _GEN_2933; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2935 = _GEN_6085 == 10'h2e2 ? _GEN_2934 : _GEN_2933; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2936 = ~io_inputBit ? 1'h0 : _GEN_2935; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2937 = _GEN_6085 == 10'h2f2 ? _GEN_2936 : _GEN_2935; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2938 = io_inputBit | _GEN_2937; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2939 = _GEN_6085 == 10'h2f2 ? _GEN_2938 : _GEN_2937; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2940 = ~io_inputBit | _GEN_2939; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2941 = _GEN_6085 == 10'h302 ? _GEN_2940 : _GEN_2939; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2942 = io_inputBit ? 1'h0 : _GEN_2941; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2943 = _GEN_6085 == 10'h302 ? _GEN_2942 : _GEN_2941; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2944 = ~io_inputBit ? 1'h0 : _GEN_2391; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2945 = i == 8'h1 ? _GEN_2944 : _GEN_2391; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2946 = io_inputBit ? 1'h0 : _GEN_2945; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2947 = i == 8'h2 ? _GEN_2946 : _GEN_2945; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2948 = io_inputBit ? 1'h0 : _GEN_2947; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2949 = i == 8'h5 ? _GEN_2948 : _GEN_2947; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2950 = ~io_inputBit ? 1'h0 : _GEN_2949; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2951 = i == 8'h9 ? _GEN_2950 : _GEN_2949; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2952 = io_inputBit ? 1'h0 : _GEN_2951; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2953 = i == 8'hb ? _GEN_2952 : _GEN_2951; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2954 = ~io_inputBit ? 1'h0 : _GEN_2953; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2955 = i == 8'h14 ? _GEN_2954 : _GEN_2953; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2956 = io_inputBit ? 1'h0 : _GEN_2955; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2957 = i == 8'h17 ? _GEN_2956 : _GEN_2955; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2958 = ~io_inputBit ? 1'h0 : _GEN_2957; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2959 = i == 8'h55 ? _GEN_2958 : _GEN_2957; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2960 = ~io_inputBit | _GEN_2959; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2961 = i == 8'h56 ? _GEN_2960 : _GEN_2959; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2962 = ~io_inputBit ? 1'h0 : _GEN_2961; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2963 = i == 8'h57 ? _GEN_2962 : _GEN_2961; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2964 = ~io_inputBit | _GEN_2963; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2965 = i == 8'h58 ? _GEN_2964 : _GEN_2963; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2966 = ~io_inputBit ? 1'h0 : _GEN_2965; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2967 = i == 8'h59 ? _GEN_2966 : _GEN_2965; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2968 = ~io_inputBit | _GEN_2967; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2969 = i == 8'h5a ? _GEN_2968 : _GEN_2967; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2970 = io_inputBit | _GEN_2969; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2971 = i == 8'h5b ? _GEN_2970 : _GEN_2969; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2972 = io_inputBit ? 1'h0 : _GEN_2971; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2973 = i == 8'h5c ? _GEN_2972 : _GEN_2971; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2974 = io_inputBit | _GEN_2973; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2975 = i == 8'h5d ? _GEN_2974 : _GEN_2973; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2976 = io_inputBit ? 1'h0 : _GEN_2975; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2977 = i == 8'h5e ? _GEN_2976 : _GEN_2975; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2978 = io_inputBit | _GEN_2977; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2979 = i == 8'h5f ? _GEN_2978 : _GEN_2977; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2980 = io_inputBit ? 1'h0 : _GEN_2979; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2981 = i == 8'h60 ? _GEN_2980 : _GEN_2979; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2982 = ~io_inputBit ? 1'h0 : _GEN_2981; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2983 = i == 8'hac ? _GEN_2982 : _GEN_2981; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2984 = ~io_inputBit | _GEN_2983; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2985 = i == 8'hae ? _GEN_2984 : _GEN_2983; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2986 = ~io_inputBit ? 1'h0 : _GEN_2985; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2987 = i == 8'hb0 ? _GEN_2986 : _GEN_2985; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2988 = ~io_inputBit | _GEN_2987; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2989 = i == 8'hb2 ? _GEN_2988 : _GEN_2987; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2990 = ~io_inputBit ? 1'h0 : _GEN_2989; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2991 = i == 8'hb4 ? _GEN_2990 : _GEN_2989; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2992 = ~io_inputBit | _GEN_2991; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2993 = i == 8'hb6 ? _GEN_2992 : _GEN_2991; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2994 = ~io_inputBit ? 1'h0 : _GEN_2993; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2995 = i == 8'hb7 ? _GEN_2994 : _GEN_2993; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2996 = ~io_inputBit | _GEN_2995; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2997 = i == 8'hb9 ? _GEN_2996 : _GEN_2995; // @[lut_mem_online.scala 235:34]
  wire  _GEN_2998 = ~io_inputBit ? 1'h0 : _GEN_2997; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_2999 = i == 8'hbb ? _GEN_2998 : _GEN_2997; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3000 = ~io_inputBit | _GEN_2999; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3001 = i == 8'hbd ? _GEN_3000 : _GEN_2999; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3002 = ~io_inputBit ? 1'h0 : _GEN_3001; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3003 = i == 8'hbf ? _GEN_3002 : _GEN_3001; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3004 = ~io_inputBit | _GEN_3003; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3005 = i == 8'hc1 ? _GEN_3004 : _GEN_3003; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3006 = ~io_inputBit ? 1'h0 : _GEN_3005; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3007 = _GEN_6084 == 9'h15a ? _GEN_3006 : _GEN_3005; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3008 = io_inputBit | _GEN_3007; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3009 = _GEN_6084 == 9'h15a ? _GEN_3008 : _GEN_3007; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3010 = ~io_inputBit | _GEN_3009; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3011 = _GEN_6084 == 9'h15e ? _GEN_3010 : _GEN_3009; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3012 = io_inputBit ? 1'h0 : _GEN_3011; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3013 = _GEN_6084 == 9'h15e ? _GEN_3012 : _GEN_3011; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3014 = ~io_inputBit ? 1'h0 : _GEN_3013; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3015 = _GEN_6084 == 9'h162 ? _GEN_3014 : _GEN_3013; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3016 = io_inputBit | _GEN_3015; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3017 = _GEN_6084 == 9'h162 ? _GEN_3016 : _GEN_3015; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3018 = ~io_inputBit | _GEN_3017; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3019 = _GEN_6084 == 9'h166 ? _GEN_3018 : _GEN_3017; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3020 = io_inputBit ? 1'h0 : _GEN_3019; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3021 = _GEN_6084 == 9'h166 ? _GEN_3020 : _GEN_3019; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3022 = ~io_inputBit ? 1'h0 : _GEN_3021; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3023 = _GEN_6084 == 9'h16a ? _GEN_3022 : _GEN_3021; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3024 = io_inputBit | _GEN_3023; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3025 = _GEN_6084 == 9'h16a ? _GEN_3024 : _GEN_3023; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3026 = ~io_inputBit | _GEN_3025; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3027 = _GEN_6084 == 9'h16e ? _GEN_3026 : _GEN_3025; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3028 = io_inputBit ? 1'h0 : _GEN_3027; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3029 = _GEN_6084 == 9'h16e ? _GEN_3028 : _GEN_3027; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3030 = ~io_inputBit ? 1'h0 : _GEN_3029; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3031 = _GEN_6084 == 9'h170 ? _GEN_3030 : _GEN_3029; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3032 = ~io_inputBit | _GEN_3031; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3033 = _GEN_6084 == 9'h174 ? _GEN_3032 : _GEN_3031; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3034 = ~io_inputBit ? 1'h0 : _GEN_3033; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3035 = _GEN_6084 == 9'h178 ? _GEN_3034 : _GEN_3033; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3036 = ~io_inputBit | _GEN_3035; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3037 = _GEN_6084 == 9'h17c ? _GEN_3036 : _GEN_3035; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3038 = ~io_inputBit ? 1'h0 : _GEN_3037; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3039 = _GEN_6084 == 9'h180 ? _GEN_3038 : _GEN_3037; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3040 = ~io_inputBit | _GEN_3039; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3041 = _GEN_6084 == 9'h184 ? _GEN_3040 : _GEN_3039; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3042 = ~io_inputBit ? 1'h0 : _GEN_3041; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3043 = _GEN_6085 == 10'h2e2 ? _GEN_3042 : _GEN_3041; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3044 = io_inputBit | _GEN_3043; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3045 = _GEN_6085 == 10'h2e2 ? _GEN_3044 : _GEN_3043; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3046 = ~io_inputBit | _GEN_3045; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3047 = _GEN_6085 == 10'h2ea ? _GEN_3046 : _GEN_3045; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3048 = io_inputBit ? 1'h0 : _GEN_3047; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3049 = _GEN_6085 == 10'h2ea ? _GEN_3048 : _GEN_3047; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3050 = ~io_inputBit ? 1'h0 : _GEN_3049; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3051 = _GEN_6085 == 10'h2f2 ? _GEN_3050 : _GEN_3049; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3052 = io_inputBit | _GEN_3051; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3053 = _GEN_6085 == 10'h2f2 ? _GEN_3052 : _GEN_3051; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3054 = ~io_inputBit | _GEN_3053; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3055 = _GEN_6085 == 10'h2fa ? _GEN_3054 : _GEN_3053; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3056 = io_inputBit ? 1'h0 : _GEN_3055; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3057 = _GEN_6085 == 10'h2fa ? _GEN_3056 : _GEN_3055; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3058 = ~io_inputBit ? 1'h0 : _GEN_3057; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3059 = _GEN_6085 == 10'h302 ? _GEN_3058 : _GEN_3057; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3060 = io_inputBit | _GEN_3059; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3061 = _GEN_6085 == 10'h302 ? _GEN_3060 : _GEN_3059; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3062 = ~io_inputBit | _GEN_3061; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3063 = _GEN_6085 == 10'h30a ? _GEN_3062 : _GEN_3061; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3064 = io_inputBit ? 1'h0 : _GEN_3063; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3065 = _GEN_6085 == 10'h30a ? _GEN_3064 : _GEN_3063; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3066 = ~io_inputBit ? 1'h0 : _GEN_2429; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3067 = i == 8'h1 ? _GEN_3066 : _GEN_2429; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3068 = io_inputBit ? 1'h0 : _GEN_3067; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3069 = i == 8'h2 ? _GEN_3068 : _GEN_3067; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3070 = io_inputBit ? 1'h0 : _GEN_3069; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3071 = i == 8'h5 ? _GEN_3070 : _GEN_3069; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3072 = ~io_inputBit ? 1'h0 : _GEN_3071; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3073 = i == 8'h9 ? _GEN_3072 : _GEN_3071; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3074 = io_inputBit ? 1'h0 : _GEN_3073; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3075 = i == 8'hb ? _GEN_3074 : _GEN_3073; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3076 = ~io_inputBit ? 1'h0 : _GEN_3075; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3077 = i == 8'h14 ? _GEN_3076 : _GEN_3075; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3078 = io_inputBit ? 1'h0 : _GEN_3077; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3079 = i == 8'h17 ? _GEN_3078 : _GEN_3077; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3080 = ~io_inputBit ? 1'h0 : _GEN_3079; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3081 = i == 8'hab ? _GEN_3080 : _GEN_3079; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3082 = ~io_inputBit | _GEN_3081; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3083 = i == 8'hac ? _GEN_3082 : _GEN_3081; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3084 = ~io_inputBit ? 1'h0 : _GEN_3083; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3085 = i == 8'had ? _GEN_3084 : _GEN_3083; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3086 = ~io_inputBit | _GEN_3085; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3087 = i == 8'hae ? _GEN_3086 : _GEN_3085; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3088 = ~io_inputBit ? 1'h0 : _GEN_3087; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3089 = i == 8'haf ? _GEN_3088 : _GEN_3087; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3090 = ~io_inputBit | _GEN_3089; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3091 = i == 8'hb0 ? _GEN_3090 : _GEN_3089; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3092 = ~io_inputBit ? 1'h0 : _GEN_3091; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3093 = i == 8'hb1 ? _GEN_3092 : _GEN_3091; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3094 = ~io_inputBit | _GEN_3093; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3095 = i == 8'hb2 ? _GEN_3094 : _GEN_3093; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3096 = ~io_inputBit ? 1'h0 : _GEN_3095; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3097 = i == 8'hb3 ? _GEN_3096 : _GEN_3095; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3098 = ~io_inputBit | _GEN_3097; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3099 = i == 8'hb4 ? _GEN_3098 : _GEN_3097; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3100 = ~io_inputBit ? 1'h0 : _GEN_3099; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3101 = i == 8'hb5 ? _GEN_3100 : _GEN_3099; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3102 = ~io_inputBit | _GEN_3101; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3103 = i == 8'hb6 ? _GEN_3102 : _GEN_3101; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3104 = ~io_inputBit ? 1'h0 : _GEN_3103; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3105 = i == 8'hb7 ? _GEN_3104 : _GEN_3103; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3106 = ~io_inputBit | _GEN_3105; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3107 = i == 8'hb8 ? _GEN_3106 : _GEN_3105; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3108 = ~io_inputBit ? 1'h0 : _GEN_3107; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3109 = i == 8'hb9 ? _GEN_3108 : _GEN_3107; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3110 = ~io_inputBit | _GEN_3109; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3111 = i == 8'hba ? _GEN_3110 : _GEN_3109; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3112 = ~io_inputBit ? 1'h0 : _GEN_3111; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3113 = i == 8'hbb ? _GEN_3112 : _GEN_3111; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3114 = ~io_inputBit | _GEN_3113; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3115 = i == 8'hbc ? _GEN_3114 : _GEN_3113; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3116 = ~io_inputBit ? 1'h0 : _GEN_3115; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3117 = i == 8'hbd ? _GEN_3116 : _GEN_3115; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3118 = ~io_inputBit | _GEN_3117; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3119 = i == 8'hbe ? _GEN_3118 : _GEN_3117; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3120 = ~io_inputBit ? 1'h0 : _GEN_3119; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3121 = i == 8'hbf ? _GEN_3120 : _GEN_3119; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3122 = ~io_inputBit | _GEN_3121; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3123 = i == 8'hc0 ? _GEN_3122 : _GEN_3121; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3124 = ~io_inputBit ? 1'h0 : _GEN_3123; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3125 = i == 8'hc1 ? _GEN_3124 : _GEN_3123; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3126 = ~io_inputBit | _GEN_3125; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3127 = i == 8'hc2 ? _GEN_3126 : _GEN_3125; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3128 = ~io_inputBit ? 1'h0 : _GEN_3127; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3129 = _GEN_6084 == 9'h158 ? _GEN_3128 : _GEN_3127; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3130 = io_inputBit | _GEN_3129; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3131 = _GEN_6084 == 9'h158 ? _GEN_3130 : _GEN_3129; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3132 = ~io_inputBit | _GEN_3131; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3133 = _GEN_6084 == 9'h15a ? _GEN_3132 : _GEN_3131; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3134 = io_inputBit ? 1'h0 : _GEN_3133; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3135 = _GEN_6084 == 9'h15a ? _GEN_3134 : _GEN_3133; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3136 = ~io_inputBit ? 1'h0 : _GEN_3135; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3137 = _GEN_6084 == 9'h15c ? _GEN_3136 : _GEN_3135; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3138 = io_inputBit | _GEN_3137; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3139 = _GEN_6084 == 9'h15c ? _GEN_3138 : _GEN_3137; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3140 = ~io_inputBit | _GEN_3139; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3141 = _GEN_6084 == 9'h15e ? _GEN_3140 : _GEN_3139; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3142 = io_inputBit ? 1'h0 : _GEN_3141; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3143 = _GEN_6084 == 9'h15e ? _GEN_3142 : _GEN_3141; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3144 = ~io_inputBit ? 1'h0 : _GEN_3143; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3145 = _GEN_6084 == 9'h160 ? _GEN_3144 : _GEN_3143; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3146 = io_inputBit | _GEN_3145; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3147 = _GEN_6084 == 9'h160 ? _GEN_3146 : _GEN_3145; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3148 = ~io_inputBit | _GEN_3147; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3149 = _GEN_6084 == 9'h162 ? _GEN_3148 : _GEN_3147; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3150 = io_inputBit ? 1'h0 : _GEN_3149; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3151 = _GEN_6084 == 9'h162 ? _GEN_3150 : _GEN_3149; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3152 = ~io_inputBit ? 1'h0 : _GEN_3151; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3153 = _GEN_6084 == 9'h164 ? _GEN_3152 : _GEN_3151; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3154 = io_inputBit | _GEN_3153; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3155 = _GEN_6084 == 9'h164 ? _GEN_3154 : _GEN_3153; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3156 = ~io_inputBit | _GEN_3155; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3157 = _GEN_6084 == 9'h166 ? _GEN_3156 : _GEN_3155; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3158 = io_inputBit ? 1'h0 : _GEN_3157; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3159 = _GEN_6084 == 9'h166 ? _GEN_3158 : _GEN_3157; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3160 = ~io_inputBit ? 1'h0 : _GEN_3159; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3161 = _GEN_6084 == 9'h168 ? _GEN_3160 : _GEN_3159; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3162 = io_inputBit | _GEN_3161; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3163 = _GEN_6084 == 9'h168 ? _GEN_3162 : _GEN_3161; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3164 = ~io_inputBit | _GEN_3163; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3165 = _GEN_6084 == 9'h16a ? _GEN_3164 : _GEN_3163; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3166 = io_inputBit ? 1'h0 : _GEN_3165; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3167 = _GEN_6084 == 9'h16a ? _GEN_3166 : _GEN_3165; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3168 = ~io_inputBit ? 1'h0 : _GEN_3167; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3169 = _GEN_6084 == 9'h16c ? _GEN_3168 : _GEN_3167; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3170 = io_inputBit | _GEN_3169; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3171 = _GEN_6084 == 9'h16c ? _GEN_3170 : _GEN_3169; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3172 = ~io_inputBit | _GEN_3171; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3173 = _GEN_6084 == 9'h16e ? _GEN_3172 : _GEN_3171; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3174 = io_inputBit ? 1'h0 : _GEN_3173; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3175 = _GEN_6084 == 9'h16e ? _GEN_3174 : _GEN_3173; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3176 = ~io_inputBit ? 1'h0 : _GEN_3175; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3177 = _GEN_6084 == 9'h170 ? _GEN_3176 : _GEN_3175; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3178 = ~io_inputBit | _GEN_3177; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3179 = _GEN_6084 == 9'h172 ? _GEN_3178 : _GEN_3177; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3180 = ~io_inputBit ? 1'h0 : _GEN_3179; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3181 = _GEN_6084 == 9'h174 ? _GEN_3180 : _GEN_3179; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3182 = ~io_inputBit | _GEN_3181; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3183 = _GEN_6084 == 9'h176 ? _GEN_3182 : _GEN_3181; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3184 = ~io_inputBit ? 1'h0 : _GEN_3183; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3185 = _GEN_6084 == 9'h178 ? _GEN_3184 : _GEN_3183; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3186 = ~io_inputBit | _GEN_3185; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3187 = _GEN_6084 == 9'h17a ? _GEN_3186 : _GEN_3185; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3188 = ~io_inputBit ? 1'h0 : _GEN_3187; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3189 = _GEN_6084 == 9'h17c ? _GEN_3188 : _GEN_3187; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3190 = ~io_inputBit | _GEN_3189; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3191 = _GEN_6084 == 9'h17e ? _GEN_3190 : _GEN_3189; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3192 = ~io_inputBit ? 1'h0 : _GEN_3191; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3193 = _GEN_6084 == 9'h180 ? _GEN_3192 : _GEN_3191; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3194 = ~io_inputBit | _GEN_3193; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3195 = _GEN_6084 == 9'h182 ? _GEN_3194 : _GEN_3193; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3196 = ~io_inputBit ? 1'h0 : _GEN_3195; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3197 = _GEN_6084 == 9'h184 ? _GEN_3196 : _GEN_3195; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3198 = ~io_inputBit | _GEN_3197; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3199 = _GEN_6084 == 9'h186 ? _GEN_3198 : _GEN_3197; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3200 = ~io_inputBit ? 1'h0 : _GEN_3199; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3201 = _GEN_6085 == 10'h2e2 ? _GEN_3200 : _GEN_3199; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3202 = io_inputBit | _GEN_3201; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3203 = _GEN_6085 == 10'h2e2 ? _GEN_3202 : _GEN_3201; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3204 = ~io_inputBit | _GEN_3203; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3205 = _GEN_6085 == 10'h2e6 ? _GEN_3204 : _GEN_3203; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3206 = io_inputBit ? 1'h0 : _GEN_3205; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3207 = _GEN_6085 == 10'h2e6 ? _GEN_3206 : _GEN_3205; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3208 = ~io_inputBit ? 1'h0 : _GEN_3207; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3209 = _GEN_6085 == 10'h2ea ? _GEN_3208 : _GEN_3207; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3210 = io_inputBit | _GEN_3209; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3211 = _GEN_6085 == 10'h2ea ? _GEN_3210 : _GEN_3209; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3212 = ~io_inputBit | _GEN_3211; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3213 = _GEN_6085 == 10'h2ee ? _GEN_3212 : _GEN_3211; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3214 = io_inputBit ? 1'h0 : _GEN_3213; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3215 = _GEN_6085 == 10'h2ee ? _GEN_3214 : _GEN_3213; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3216 = ~io_inputBit ? 1'h0 : _GEN_3215; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3217 = _GEN_6085 == 10'h2f2 ? _GEN_3216 : _GEN_3215; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3218 = io_inputBit | _GEN_3217; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3219 = _GEN_6085 == 10'h2f2 ? _GEN_3218 : _GEN_3217; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3220 = ~io_inputBit | _GEN_3219; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3221 = _GEN_6085 == 10'h2f6 ? _GEN_3220 : _GEN_3219; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3222 = io_inputBit ? 1'h0 : _GEN_3221; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3223 = _GEN_6085 == 10'h2f6 ? _GEN_3222 : _GEN_3221; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3224 = ~io_inputBit ? 1'h0 : _GEN_3223; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3225 = _GEN_6085 == 10'h2fa ? _GEN_3224 : _GEN_3223; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3226 = io_inputBit | _GEN_3225; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3227 = _GEN_6085 == 10'h2fa ? _GEN_3226 : _GEN_3225; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3228 = ~io_inputBit | _GEN_3227; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3229 = _GEN_6085 == 10'h2fe ? _GEN_3228 : _GEN_3227; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3230 = io_inputBit ? 1'h0 : _GEN_3229; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3231 = _GEN_6085 == 10'h2fe ? _GEN_3230 : _GEN_3229; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3232 = ~io_inputBit ? 1'h0 : _GEN_3231; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3233 = _GEN_6085 == 10'h302 ? _GEN_3232 : _GEN_3231; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3234 = io_inputBit | _GEN_3233; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3235 = _GEN_6085 == 10'h302 ? _GEN_3234 : _GEN_3233; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3236 = ~io_inputBit | _GEN_3235; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3237 = _GEN_6085 == 10'h306 ? _GEN_3236 : _GEN_3235; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3238 = io_inputBit ? 1'h0 : _GEN_3237; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3239 = _GEN_6085 == 10'h306 ? _GEN_3238 : _GEN_3237; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3240 = ~io_inputBit ? 1'h0 : _GEN_3239; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3241 = _GEN_6085 == 10'h30a ? _GEN_3240 : _GEN_3239; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3242 = io_inputBit | _GEN_3241; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3243 = _GEN_6085 == 10'h30a ? _GEN_3242 : _GEN_3241; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3244 = ~io_inputBit | _GEN_3243; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3245 = _GEN_6085 == 10'h30e ? _GEN_3244 : _GEN_3243; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3246 = io_inputBit ? 1'h0 : _GEN_3245; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3247 = _GEN_6085 == 10'h30e ? _GEN_3246 : _GEN_3245; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3248 = ~io_inputBit ? 1'h0 : _GEN_2499; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3249 = i == 8'h1 ? _GEN_3248 : _GEN_2499; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3250 = io_inputBit ? 1'h0 : _GEN_3249; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3251 = i == 8'h2 ? _GEN_3250 : _GEN_3249; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3252 = io_inputBit ? 1'h0 : _GEN_3251; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3253 = i == 8'h5 ? _GEN_3252 : _GEN_3251; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3254 = ~io_inputBit ? 1'h0 : _GEN_3253; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3255 = i == 8'h9 ? _GEN_3254 : _GEN_3253; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3256 = io_inputBit ? 1'h0 : _GEN_3255; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3257 = i == 8'hb ? _GEN_3256 : _GEN_3255; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3258 = ~io_inputBit ? 1'h0 : _GEN_3257; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3259 = i == 8'h14 ? _GEN_3258 : _GEN_3257; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3260 = io_inputBit ? 1'h0 : _GEN_3259; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3261 = i == 8'h30 ? _GEN_3260 : _GEN_3259; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3262 = io_inputBit ? 1'h0 : _GEN_3261; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3263 = i == 8'h61 ? _GEN_3262 : _GEN_3261; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3264 = io_inputBit ? 1'h0 : _GEN_3263; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3265 = i == 8'hc3 ? _GEN_3264 : _GEN_3263; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3266 = ~io_inputBit ? 1'h0 : _GEN_3265; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3267 = _GEN_6084 == 9'h157 ? _GEN_3266 : _GEN_3265; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3268 = io_inputBit | _GEN_3267; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3269 = _GEN_6084 == 9'h157 ? _GEN_3268 : _GEN_3267; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3270 = ~io_inputBit | _GEN_3269; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3271 = _GEN_6084 == 9'h158 ? _GEN_3270 : _GEN_3269; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3272 = io_inputBit ? 1'h0 : _GEN_3271; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3273 = _GEN_6084 == 9'h158 ? _GEN_3272 : _GEN_3271; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3274 = ~io_inputBit ? 1'h0 : _GEN_3273; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3275 = _GEN_6084 == 9'h159 ? _GEN_3274 : _GEN_3273; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3276 = io_inputBit | _GEN_3275; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3277 = _GEN_6084 == 9'h159 ? _GEN_3276 : _GEN_3275; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3278 = ~io_inputBit | _GEN_3277; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3279 = _GEN_6084 == 9'h15a ? _GEN_3278 : _GEN_3277; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3280 = io_inputBit ? 1'h0 : _GEN_3279; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3281 = _GEN_6084 == 9'h15a ? _GEN_3280 : _GEN_3279; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3282 = ~io_inputBit ? 1'h0 : _GEN_3281; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3283 = _GEN_6084 == 9'h15b ? _GEN_3282 : _GEN_3281; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3284 = io_inputBit | _GEN_3283; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3285 = _GEN_6084 == 9'h15b ? _GEN_3284 : _GEN_3283; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3286 = ~io_inputBit | _GEN_3285; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3287 = _GEN_6084 == 9'h15c ? _GEN_3286 : _GEN_3285; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3288 = io_inputBit ? 1'h0 : _GEN_3287; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3289 = _GEN_6084 == 9'h15c ? _GEN_3288 : _GEN_3287; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3290 = ~io_inputBit ? 1'h0 : _GEN_3289; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3291 = _GEN_6084 == 9'h15d ? _GEN_3290 : _GEN_3289; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3292 = io_inputBit | _GEN_3291; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3293 = _GEN_6084 == 9'h15d ? _GEN_3292 : _GEN_3291; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3294 = ~io_inputBit | _GEN_3293; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3295 = _GEN_6084 == 9'h15e ? _GEN_3294 : _GEN_3293; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3296 = io_inputBit ? 1'h0 : _GEN_3295; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3297 = _GEN_6084 == 9'h15e ? _GEN_3296 : _GEN_3295; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3298 = ~io_inputBit ? 1'h0 : _GEN_3297; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3299 = _GEN_6084 == 9'h15f ? _GEN_3298 : _GEN_3297; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3300 = io_inputBit | _GEN_3299; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3301 = _GEN_6084 == 9'h15f ? _GEN_3300 : _GEN_3299; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3302 = ~io_inputBit | _GEN_3301; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3303 = _GEN_6084 == 9'h160 ? _GEN_3302 : _GEN_3301; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3304 = io_inputBit ? 1'h0 : _GEN_3303; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3305 = _GEN_6084 == 9'h160 ? _GEN_3304 : _GEN_3303; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3306 = ~io_inputBit ? 1'h0 : _GEN_3305; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3307 = _GEN_6084 == 9'h161 ? _GEN_3306 : _GEN_3305; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3308 = io_inputBit | _GEN_3307; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3309 = _GEN_6084 == 9'h161 ? _GEN_3308 : _GEN_3307; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3310 = ~io_inputBit | _GEN_3309; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3311 = _GEN_6084 == 9'h162 ? _GEN_3310 : _GEN_3309; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3312 = io_inputBit ? 1'h0 : _GEN_3311; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3313 = _GEN_6084 == 9'h162 ? _GEN_3312 : _GEN_3311; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3314 = ~io_inputBit ? 1'h0 : _GEN_3313; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3315 = _GEN_6084 == 9'h163 ? _GEN_3314 : _GEN_3313; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3316 = io_inputBit | _GEN_3315; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3317 = _GEN_6084 == 9'h163 ? _GEN_3316 : _GEN_3315; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3318 = ~io_inputBit | _GEN_3317; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3319 = _GEN_6084 == 9'h164 ? _GEN_3318 : _GEN_3317; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3320 = io_inputBit ? 1'h0 : _GEN_3319; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3321 = _GEN_6084 == 9'h164 ? _GEN_3320 : _GEN_3319; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3322 = ~io_inputBit ? 1'h0 : _GEN_3321; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3323 = _GEN_6084 == 9'h165 ? _GEN_3322 : _GEN_3321; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3324 = io_inputBit | _GEN_3323; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3325 = _GEN_6084 == 9'h165 ? _GEN_3324 : _GEN_3323; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3326 = ~io_inputBit | _GEN_3325; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3327 = _GEN_6084 == 9'h166 ? _GEN_3326 : _GEN_3325; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3328 = io_inputBit ? 1'h0 : _GEN_3327; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3329 = _GEN_6084 == 9'h166 ? _GEN_3328 : _GEN_3327; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3330 = ~io_inputBit ? 1'h0 : _GEN_3329; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3331 = _GEN_6084 == 9'h167 ? _GEN_3330 : _GEN_3329; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3332 = io_inputBit | _GEN_3331; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3333 = _GEN_6084 == 9'h167 ? _GEN_3332 : _GEN_3331; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3334 = ~io_inputBit | _GEN_3333; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3335 = _GEN_6084 == 9'h168 ? _GEN_3334 : _GEN_3333; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3336 = io_inputBit ? 1'h0 : _GEN_3335; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3337 = _GEN_6084 == 9'h168 ? _GEN_3336 : _GEN_3335; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3338 = ~io_inputBit ? 1'h0 : _GEN_3337; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3339 = _GEN_6084 == 9'h169 ? _GEN_3338 : _GEN_3337; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3340 = io_inputBit | _GEN_3339; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3341 = _GEN_6084 == 9'h169 ? _GEN_3340 : _GEN_3339; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3342 = ~io_inputBit | _GEN_3341; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3343 = _GEN_6084 == 9'h16a ? _GEN_3342 : _GEN_3341; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3344 = io_inputBit ? 1'h0 : _GEN_3343; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3345 = _GEN_6084 == 9'h16a ? _GEN_3344 : _GEN_3343; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3346 = ~io_inputBit ? 1'h0 : _GEN_3345; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3347 = _GEN_6084 == 9'h16b ? _GEN_3346 : _GEN_3345; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3348 = io_inputBit | _GEN_3347; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3349 = _GEN_6084 == 9'h16b ? _GEN_3348 : _GEN_3347; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3350 = ~io_inputBit | _GEN_3349; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3351 = _GEN_6084 == 9'h16c ? _GEN_3350 : _GEN_3349; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3352 = io_inputBit ? 1'h0 : _GEN_3351; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3353 = _GEN_6084 == 9'h16c ? _GEN_3352 : _GEN_3351; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3354 = ~io_inputBit ? 1'h0 : _GEN_3353; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3355 = _GEN_6084 == 9'h16d ? _GEN_3354 : _GEN_3353; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3356 = io_inputBit | _GEN_3355; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3357 = _GEN_6084 == 9'h16d ? _GEN_3356 : _GEN_3355; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3358 = ~io_inputBit | _GEN_3357; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3359 = _GEN_6084 == 9'h16e ? _GEN_3358 : _GEN_3357; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3360 = io_inputBit ? 1'h0 : _GEN_3359; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3361 = _GEN_6084 == 9'h16e ? _GEN_3360 : _GEN_3359; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3362 = ~io_inputBit ? 1'h0 : _GEN_3361; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3363 = _GEN_6084 == 9'h16f ? _GEN_3362 : _GEN_3361; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3364 = ~io_inputBit ? 1'h0 : _GEN_3363; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3365 = _GEN_6084 == 9'h170 ? _GEN_3364 : _GEN_3363; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3366 = ~io_inputBit | _GEN_3365; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3367 = _GEN_6084 == 9'h171 ? _GEN_3366 : _GEN_3365; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3368 = ~io_inputBit ? 1'h0 : _GEN_3367; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3369 = _GEN_6084 == 9'h172 ? _GEN_3368 : _GEN_3367; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3370 = ~io_inputBit | _GEN_3369; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3371 = _GEN_6084 == 9'h173 ? _GEN_3370 : _GEN_3369; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3372 = ~io_inputBit ? 1'h0 : _GEN_3371; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3373 = _GEN_6084 == 9'h174 ? _GEN_3372 : _GEN_3371; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3374 = ~io_inputBit | _GEN_3373; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3375 = _GEN_6084 == 9'h175 ? _GEN_3374 : _GEN_3373; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3376 = ~io_inputBit ? 1'h0 : _GEN_3375; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3377 = _GEN_6084 == 9'h176 ? _GEN_3376 : _GEN_3375; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3378 = ~io_inputBit | _GEN_3377; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3379 = _GEN_6084 == 9'h177 ? _GEN_3378 : _GEN_3377; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3380 = ~io_inputBit ? 1'h0 : _GEN_3379; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3381 = _GEN_6084 == 9'h178 ? _GEN_3380 : _GEN_3379; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3382 = ~io_inputBit | _GEN_3381; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3383 = _GEN_6084 == 9'h179 ? _GEN_3382 : _GEN_3381; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3384 = ~io_inputBit ? 1'h0 : _GEN_3383; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3385 = _GEN_6084 == 9'h17a ? _GEN_3384 : _GEN_3383; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3386 = ~io_inputBit | _GEN_3385; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3387 = _GEN_6084 == 9'h17b ? _GEN_3386 : _GEN_3385; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3388 = ~io_inputBit ? 1'h0 : _GEN_3387; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3389 = _GEN_6084 == 9'h17c ? _GEN_3388 : _GEN_3387; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3390 = ~io_inputBit | _GEN_3389; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3391 = _GEN_6084 == 9'h17d ? _GEN_3390 : _GEN_3389; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3392 = ~io_inputBit ? 1'h0 : _GEN_3391; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3393 = _GEN_6084 == 9'h17e ? _GEN_3392 : _GEN_3391; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3394 = ~io_inputBit | _GEN_3393; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3395 = _GEN_6084 == 9'h17f ? _GEN_3394 : _GEN_3393; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3396 = ~io_inputBit ? 1'h0 : _GEN_3395; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3397 = _GEN_6084 == 9'h180 ? _GEN_3396 : _GEN_3395; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3398 = ~io_inputBit | _GEN_3397; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3399 = _GEN_6084 == 9'h181 ? _GEN_3398 : _GEN_3397; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3400 = ~io_inputBit ? 1'h0 : _GEN_3399; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3401 = _GEN_6084 == 9'h182 ? _GEN_3400 : _GEN_3399; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3402 = ~io_inputBit | _GEN_3401; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3403 = _GEN_6084 == 9'h183 ? _GEN_3402 : _GEN_3401; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3404 = ~io_inputBit ? 1'h0 : _GEN_3403; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3405 = _GEN_6084 == 9'h184 ? _GEN_3404 : _GEN_3403; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3406 = ~io_inputBit | _GEN_3405; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3407 = _GEN_6084 == 9'h185 ? _GEN_3406 : _GEN_3405; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3408 = ~io_inputBit ? 1'h0 : _GEN_3407; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3409 = _GEN_6084 == 9'h186 ? _GEN_3408 : _GEN_3407; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3410 = ~io_inputBit | _GEN_3409; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3411 = _GEN_6084 == 9'h187 ? _GEN_3410 : _GEN_3409; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3412 = ~io_inputBit | _GEN_3411; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3413 = _GEN_6085 == 10'h2e0 ? _GEN_3412 : _GEN_3411; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3414 = io_inputBit ? 1'h0 : _GEN_3413; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3415 = _GEN_6085 == 10'h2e0 ? _GEN_3414 : _GEN_3413; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3416 = ~io_inputBit ? 1'h0 : _GEN_3415; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3417 = _GEN_6085 == 10'h2e2 ? _GEN_3416 : _GEN_3415; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3418 = io_inputBit | _GEN_3417; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3419 = _GEN_6085 == 10'h2e2 ? _GEN_3418 : _GEN_3417; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3420 = ~io_inputBit | _GEN_3419; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3421 = _GEN_6085 == 10'h2e4 ? _GEN_3420 : _GEN_3419; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3422 = io_inputBit ? 1'h0 : _GEN_3421; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3423 = _GEN_6085 == 10'h2e4 ? _GEN_3422 : _GEN_3421; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3424 = ~io_inputBit ? 1'h0 : _GEN_3423; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3425 = _GEN_6085 == 10'h2e6 ? _GEN_3424 : _GEN_3423; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3426 = io_inputBit | _GEN_3425; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3427 = _GEN_6085 == 10'h2e6 ? _GEN_3426 : _GEN_3425; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3428 = ~io_inputBit | _GEN_3427; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3429 = _GEN_6085 == 10'h2e8 ? _GEN_3428 : _GEN_3427; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3430 = io_inputBit ? 1'h0 : _GEN_3429; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3431 = _GEN_6085 == 10'h2e8 ? _GEN_3430 : _GEN_3429; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3432 = ~io_inputBit ? 1'h0 : _GEN_3431; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3433 = _GEN_6085 == 10'h2ea ? _GEN_3432 : _GEN_3431; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3434 = io_inputBit | _GEN_3433; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3435 = _GEN_6085 == 10'h2ea ? _GEN_3434 : _GEN_3433; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3436 = ~io_inputBit | _GEN_3435; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3437 = _GEN_6085 == 10'h2ec ? _GEN_3436 : _GEN_3435; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3438 = io_inputBit ? 1'h0 : _GEN_3437; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3439 = _GEN_6085 == 10'h2ec ? _GEN_3438 : _GEN_3437; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3440 = ~io_inputBit ? 1'h0 : _GEN_3439; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3441 = _GEN_6085 == 10'h2ee ? _GEN_3440 : _GEN_3439; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3442 = io_inputBit | _GEN_3441; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3443 = _GEN_6085 == 10'h2ee ? _GEN_3442 : _GEN_3441; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3444 = ~io_inputBit | _GEN_3443; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3445 = _GEN_6085 == 10'h2f0 ? _GEN_3444 : _GEN_3443; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3446 = io_inputBit ? 1'h0 : _GEN_3445; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3447 = _GEN_6085 == 10'h2f0 ? _GEN_3446 : _GEN_3445; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3448 = ~io_inputBit ? 1'h0 : _GEN_3447; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3449 = _GEN_6085 == 10'h2f2 ? _GEN_3448 : _GEN_3447; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3450 = io_inputBit | _GEN_3449; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3451 = _GEN_6085 == 10'h2f2 ? _GEN_3450 : _GEN_3449; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3452 = ~io_inputBit | _GEN_3451; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3453 = _GEN_6085 == 10'h2f4 ? _GEN_3452 : _GEN_3451; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3454 = io_inputBit ? 1'h0 : _GEN_3453; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3455 = _GEN_6085 == 10'h2f4 ? _GEN_3454 : _GEN_3453; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3456 = ~io_inputBit ? 1'h0 : _GEN_3455; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3457 = _GEN_6085 == 10'h2f6 ? _GEN_3456 : _GEN_3455; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3458 = io_inputBit | _GEN_3457; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3459 = _GEN_6085 == 10'h2f6 ? _GEN_3458 : _GEN_3457; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3460 = ~io_inputBit | _GEN_3459; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3461 = _GEN_6085 == 10'h2f8 ? _GEN_3460 : _GEN_3459; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3462 = io_inputBit ? 1'h0 : _GEN_3461; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3463 = _GEN_6085 == 10'h2f8 ? _GEN_3462 : _GEN_3461; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3464 = ~io_inputBit ? 1'h0 : _GEN_3463; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3465 = _GEN_6085 == 10'h2fa ? _GEN_3464 : _GEN_3463; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3466 = io_inputBit | _GEN_3465; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3467 = _GEN_6085 == 10'h2fa ? _GEN_3466 : _GEN_3465; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3468 = ~io_inputBit | _GEN_3467; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3469 = _GEN_6085 == 10'h2fc ? _GEN_3468 : _GEN_3467; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3470 = io_inputBit ? 1'h0 : _GEN_3469; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3471 = _GEN_6085 == 10'h2fc ? _GEN_3470 : _GEN_3469; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3472 = ~io_inputBit ? 1'h0 : _GEN_3471; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3473 = _GEN_6085 == 10'h2fe ? _GEN_3472 : _GEN_3471; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3474 = io_inputBit | _GEN_3473; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3475 = _GEN_6085 == 10'h2fe ? _GEN_3474 : _GEN_3473; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3476 = ~io_inputBit | _GEN_3475; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3477 = _GEN_6085 == 10'h300 ? _GEN_3476 : _GEN_3475; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3478 = io_inputBit ? 1'h0 : _GEN_3477; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3479 = _GEN_6085 == 10'h300 ? _GEN_3478 : _GEN_3477; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3480 = ~io_inputBit ? 1'h0 : _GEN_3479; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3481 = _GEN_6085 == 10'h302 ? _GEN_3480 : _GEN_3479; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3482 = io_inputBit | _GEN_3481; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3483 = _GEN_6085 == 10'h302 ? _GEN_3482 : _GEN_3481; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3484 = ~io_inputBit | _GEN_3483; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3485 = _GEN_6085 == 10'h304 ? _GEN_3484 : _GEN_3483; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3486 = io_inputBit ? 1'h0 : _GEN_3485; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3487 = _GEN_6085 == 10'h304 ? _GEN_3486 : _GEN_3485; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3488 = ~io_inputBit ? 1'h0 : _GEN_3487; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3489 = _GEN_6085 == 10'h306 ? _GEN_3488 : _GEN_3487; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3490 = io_inputBit | _GEN_3489; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3491 = _GEN_6085 == 10'h306 ? _GEN_3490 : _GEN_3489; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3492 = ~io_inputBit | _GEN_3491; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3493 = _GEN_6085 == 10'h308 ? _GEN_3492 : _GEN_3491; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3494 = io_inputBit ? 1'h0 : _GEN_3493; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3495 = _GEN_6085 == 10'h308 ? _GEN_3494 : _GEN_3493; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3496 = ~io_inputBit ? 1'h0 : _GEN_3495; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3497 = _GEN_6085 == 10'h30a ? _GEN_3496 : _GEN_3495; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3498 = io_inputBit | _GEN_3497; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3499 = _GEN_6085 == 10'h30a ? _GEN_3498 : _GEN_3497; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3500 = ~io_inputBit | _GEN_3499; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3501 = _GEN_6085 == 10'h30c ? _GEN_3500 : _GEN_3499; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3502 = io_inputBit ? 1'h0 : _GEN_3501; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3503 = _GEN_6085 == 10'h30c ? _GEN_3502 : _GEN_3501; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3504 = ~io_inputBit ? 1'h0 : _GEN_3503; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3505 = _GEN_6085 == 10'h30e ? _GEN_3504 : _GEN_3503; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3506 = io_inputBit | _GEN_3505; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3507 = _GEN_6085 == 10'h30e ? _GEN_3506 : _GEN_3505; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3508 = ~io_inputBit | _GEN_3507; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3509 = _GEN_6085 == 10'h310 ? _GEN_3508 : _GEN_3507; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3510 = io_inputBit ? 1'h0 : _GEN_3509; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3511 = _GEN_6085 == 10'h310 ? _GEN_3510 : _GEN_3509; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3512 = ~io_inputBit ? 1'h0 : _GEN_2615; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3513 = i == 8'h1 ? _GEN_3512 : _GEN_2615; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3514 = io_inputBit ? 1'h0 : _GEN_3513; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3515 = i == 8'h2 ? _GEN_3514 : _GEN_3513; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3516 = io_inputBit ? 1'h0 : _GEN_3515; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3517 = i == 8'h5 ? _GEN_3516 : _GEN_3515; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3518 = ~io_inputBit ? 1'h0 : _GEN_3517; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3519 = i == 8'h9 ? _GEN_3518 : _GEN_3517; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3520 = io_inputBit ? 1'h0 : _GEN_3519; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3521 = i == 8'hb ? _GEN_3520 : _GEN_3519; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3522 = ~io_inputBit ? 1'h0 : _GEN_3521; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3523 = i == 8'h14 ? _GEN_3522 : _GEN_3521; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3524 = io_inputBit ? 1'h0 : _GEN_3523; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3525 = i == 8'h30 ? _GEN_3524 : _GEN_3523; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3526 = io_inputBit ? 1'h0 : _GEN_3525; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3527 = i == 8'h61 ? _GEN_3526 : _GEN_3525; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3528 = ~io_inputBit | _GEN_3527; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3529 = _GEN_6084 == 9'h157 ? _GEN_3528 : _GEN_3527; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3530 = io_inputBit ? 1'h0 : _GEN_3529; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3531 = _GEN_6084 == 9'h157 ? _GEN_3530 : _GEN_3529; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3532 = ~io_inputBit | _GEN_3531; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3533 = _GEN_6084 == 9'h158 ? _GEN_3532 : _GEN_3531; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3534 = io_inputBit ? 1'h0 : _GEN_3533; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3535 = _GEN_6084 == 9'h158 ? _GEN_3534 : _GEN_3533; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3536 = ~io_inputBit | _GEN_3535; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3537 = _GEN_6084 == 9'h159 ? _GEN_3536 : _GEN_3535; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3538 = io_inputBit ? 1'h0 : _GEN_3537; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3539 = _GEN_6084 == 9'h159 ? _GEN_3538 : _GEN_3537; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3540 = ~io_inputBit | _GEN_3539; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3541 = _GEN_6084 == 9'h15a ? _GEN_3540 : _GEN_3539; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3542 = io_inputBit ? 1'h0 : _GEN_3541; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3543 = _GEN_6084 == 9'h15a ? _GEN_3542 : _GEN_3541; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3544 = ~io_inputBit | _GEN_3543; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3545 = _GEN_6084 == 9'h15b ? _GEN_3544 : _GEN_3543; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3546 = io_inputBit ? 1'h0 : _GEN_3545; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3547 = _GEN_6084 == 9'h15b ? _GEN_3546 : _GEN_3545; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3548 = ~io_inputBit | _GEN_3547; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3549 = _GEN_6084 == 9'h15c ? _GEN_3548 : _GEN_3547; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3550 = io_inputBit ? 1'h0 : _GEN_3549; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3551 = _GEN_6084 == 9'h15c ? _GEN_3550 : _GEN_3549; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3552 = ~io_inputBit | _GEN_3551; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3553 = _GEN_6084 == 9'h15d ? _GEN_3552 : _GEN_3551; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3554 = io_inputBit ? 1'h0 : _GEN_3553; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3555 = _GEN_6084 == 9'h15d ? _GEN_3554 : _GEN_3553; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3556 = ~io_inputBit | _GEN_3555; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3557 = _GEN_6084 == 9'h15e ? _GEN_3556 : _GEN_3555; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3558 = io_inputBit ? 1'h0 : _GEN_3557; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3559 = _GEN_6084 == 9'h15e ? _GEN_3558 : _GEN_3557; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3560 = ~io_inputBit | _GEN_3559; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3561 = _GEN_6084 == 9'h15f ? _GEN_3560 : _GEN_3559; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3562 = io_inputBit ? 1'h0 : _GEN_3561; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3563 = _GEN_6084 == 9'h15f ? _GEN_3562 : _GEN_3561; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3564 = ~io_inputBit | _GEN_3563; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3565 = _GEN_6084 == 9'h160 ? _GEN_3564 : _GEN_3563; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3566 = io_inputBit ? 1'h0 : _GEN_3565; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3567 = _GEN_6084 == 9'h160 ? _GEN_3566 : _GEN_3565; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3568 = ~io_inputBit | _GEN_3567; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3569 = _GEN_6084 == 9'h161 ? _GEN_3568 : _GEN_3567; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3570 = io_inputBit ? 1'h0 : _GEN_3569; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3571 = _GEN_6084 == 9'h161 ? _GEN_3570 : _GEN_3569; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3572 = ~io_inputBit | _GEN_3571; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3573 = _GEN_6084 == 9'h162 ? _GEN_3572 : _GEN_3571; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3574 = io_inputBit ? 1'h0 : _GEN_3573; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3575 = _GEN_6084 == 9'h162 ? _GEN_3574 : _GEN_3573; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3576 = ~io_inputBit | _GEN_3575; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3577 = _GEN_6084 == 9'h163 ? _GEN_3576 : _GEN_3575; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3578 = io_inputBit ? 1'h0 : _GEN_3577; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3579 = _GEN_6084 == 9'h163 ? _GEN_3578 : _GEN_3577; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3580 = ~io_inputBit | _GEN_3579; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3581 = _GEN_6084 == 9'h164 ? _GEN_3580 : _GEN_3579; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3582 = io_inputBit ? 1'h0 : _GEN_3581; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3583 = _GEN_6084 == 9'h164 ? _GEN_3582 : _GEN_3581; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3584 = ~io_inputBit | _GEN_3583; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3585 = _GEN_6084 == 9'h165 ? _GEN_3584 : _GEN_3583; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3586 = io_inputBit ? 1'h0 : _GEN_3585; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3587 = _GEN_6084 == 9'h165 ? _GEN_3586 : _GEN_3585; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3588 = ~io_inputBit | _GEN_3587; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3589 = _GEN_6084 == 9'h166 ? _GEN_3588 : _GEN_3587; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3590 = io_inputBit ? 1'h0 : _GEN_3589; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3591 = _GEN_6084 == 9'h166 ? _GEN_3590 : _GEN_3589; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3592 = ~io_inputBit | _GEN_3591; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3593 = _GEN_6084 == 9'h167 ? _GEN_3592 : _GEN_3591; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3594 = io_inputBit ? 1'h0 : _GEN_3593; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3595 = _GEN_6084 == 9'h167 ? _GEN_3594 : _GEN_3593; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3596 = ~io_inputBit | _GEN_3595; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3597 = _GEN_6084 == 9'h168 ? _GEN_3596 : _GEN_3595; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3598 = io_inputBit ? 1'h0 : _GEN_3597; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3599 = _GEN_6084 == 9'h168 ? _GEN_3598 : _GEN_3597; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3600 = ~io_inputBit | _GEN_3599; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3601 = _GEN_6084 == 9'h169 ? _GEN_3600 : _GEN_3599; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3602 = io_inputBit ? 1'h0 : _GEN_3601; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3603 = _GEN_6084 == 9'h169 ? _GEN_3602 : _GEN_3601; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3604 = ~io_inputBit | _GEN_3603; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3605 = _GEN_6084 == 9'h16a ? _GEN_3604 : _GEN_3603; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3606 = io_inputBit ? 1'h0 : _GEN_3605; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3607 = _GEN_6084 == 9'h16a ? _GEN_3606 : _GEN_3605; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3608 = ~io_inputBit | _GEN_3607; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3609 = _GEN_6084 == 9'h16b ? _GEN_3608 : _GEN_3607; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3610 = io_inputBit ? 1'h0 : _GEN_3609; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3611 = _GEN_6084 == 9'h16b ? _GEN_3610 : _GEN_3609; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3612 = ~io_inputBit | _GEN_3611; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3613 = _GEN_6084 == 9'h16c ? _GEN_3612 : _GEN_3611; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3614 = io_inputBit ? 1'h0 : _GEN_3613; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3615 = _GEN_6084 == 9'h16c ? _GEN_3614 : _GEN_3613; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3616 = ~io_inputBit | _GEN_3615; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3617 = _GEN_6084 == 9'h16d ? _GEN_3616 : _GEN_3615; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3618 = io_inputBit ? 1'h0 : _GEN_3617; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3619 = _GEN_6084 == 9'h16d ? _GEN_3618 : _GEN_3617; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3620 = ~io_inputBit | _GEN_3619; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3621 = _GEN_6084 == 9'h16e ? _GEN_3620 : _GEN_3619; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3622 = io_inputBit ? 1'h0 : _GEN_3621; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3623 = _GEN_6084 == 9'h16e ? _GEN_3622 : _GEN_3621; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3624 = ~io_inputBit | _GEN_3623; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3625 = _GEN_6084 == 9'h16f ? _GEN_3624 : _GEN_3623; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3626 = io_inputBit ? 1'h0 : _GEN_3625; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3627 = _GEN_6084 == 9'h188 ? _GEN_3626 : _GEN_3625; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3628 = ~io_inputBit ? 1'h0 : _GEN_3627; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3629 = _GEN_6085 == 10'h2e0 ? _GEN_3628 : _GEN_3627; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3630 = io_inputBit | _GEN_3629; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3631 = _GEN_6085 == 10'h2e0 ? _GEN_3630 : _GEN_3629; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3632 = ~io_inputBit | _GEN_3631; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3633 = _GEN_6085 == 10'h2e1 ? _GEN_3632 : _GEN_3631; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3634 = io_inputBit ? 1'h0 : _GEN_3633; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3635 = _GEN_6085 == 10'h2e1 ? _GEN_3634 : _GEN_3633; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3636 = ~io_inputBit ? 1'h0 : _GEN_3635; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3637 = _GEN_6085 == 10'h2e2 ? _GEN_3636 : _GEN_3635; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3638 = io_inputBit | _GEN_3637; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3639 = _GEN_6085 == 10'h2e2 ? _GEN_3638 : _GEN_3637; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3640 = ~io_inputBit | _GEN_3639; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3641 = _GEN_6085 == 10'h2e3 ? _GEN_3640 : _GEN_3639; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3642 = io_inputBit ? 1'h0 : _GEN_3641; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3643 = _GEN_6085 == 10'h2e3 ? _GEN_3642 : _GEN_3641; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3644 = ~io_inputBit ? 1'h0 : _GEN_3643; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3645 = _GEN_6085 == 10'h2e4 ? _GEN_3644 : _GEN_3643; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3646 = io_inputBit | _GEN_3645; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3647 = _GEN_6085 == 10'h2e4 ? _GEN_3646 : _GEN_3645; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3648 = ~io_inputBit | _GEN_3647; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3649 = _GEN_6085 == 10'h2e5 ? _GEN_3648 : _GEN_3647; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3650 = io_inputBit ? 1'h0 : _GEN_3649; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3651 = _GEN_6085 == 10'h2e5 ? _GEN_3650 : _GEN_3649; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3652 = ~io_inputBit ? 1'h0 : _GEN_3651; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3653 = _GEN_6085 == 10'h2e6 ? _GEN_3652 : _GEN_3651; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3654 = io_inputBit | _GEN_3653; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3655 = _GEN_6085 == 10'h2e6 ? _GEN_3654 : _GEN_3653; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3656 = ~io_inputBit | _GEN_3655; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3657 = _GEN_6085 == 10'h2e7 ? _GEN_3656 : _GEN_3655; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3658 = io_inputBit ? 1'h0 : _GEN_3657; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3659 = _GEN_6085 == 10'h2e7 ? _GEN_3658 : _GEN_3657; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3660 = ~io_inputBit ? 1'h0 : _GEN_3659; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3661 = _GEN_6085 == 10'h2e8 ? _GEN_3660 : _GEN_3659; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3662 = io_inputBit | _GEN_3661; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3663 = _GEN_6085 == 10'h2e8 ? _GEN_3662 : _GEN_3661; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3664 = ~io_inputBit | _GEN_3663; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3665 = _GEN_6085 == 10'h2e9 ? _GEN_3664 : _GEN_3663; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3666 = io_inputBit ? 1'h0 : _GEN_3665; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3667 = _GEN_6085 == 10'h2e9 ? _GEN_3666 : _GEN_3665; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3668 = ~io_inputBit ? 1'h0 : _GEN_3667; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3669 = _GEN_6085 == 10'h2ea ? _GEN_3668 : _GEN_3667; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3670 = io_inputBit | _GEN_3669; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3671 = _GEN_6085 == 10'h2ea ? _GEN_3670 : _GEN_3669; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3672 = ~io_inputBit | _GEN_3671; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3673 = _GEN_6085 == 10'h2eb ? _GEN_3672 : _GEN_3671; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3674 = io_inputBit ? 1'h0 : _GEN_3673; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3675 = _GEN_6085 == 10'h2eb ? _GEN_3674 : _GEN_3673; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3676 = ~io_inputBit ? 1'h0 : _GEN_3675; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3677 = _GEN_6085 == 10'h2ec ? _GEN_3676 : _GEN_3675; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3678 = io_inputBit | _GEN_3677; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3679 = _GEN_6085 == 10'h2ec ? _GEN_3678 : _GEN_3677; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3680 = ~io_inputBit | _GEN_3679; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3681 = _GEN_6085 == 10'h2ed ? _GEN_3680 : _GEN_3679; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3682 = io_inputBit ? 1'h0 : _GEN_3681; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3683 = _GEN_6085 == 10'h2ed ? _GEN_3682 : _GEN_3681; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3684 = ~io_inputBit ? 1'h0 : _GEN_3683; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3685 = _GEN_6085 == 10'h2ee ? _GEN_3684 : _GEN_3683; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3686 = io_inputBit | _GEN_3685; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3687 = _GEN_6085 == 10'h2ee ? _GEN_3686 : _GEN_3685; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3688 = ~io_inputBit | _GEN_3687; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3689 = _GEN_6085 == 10'h2ef ? _GEN_3688 : _GEN_3687; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3690 = io_inputBit ? 1'h0 : _GEN_3689; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3691 = _GEN_6085 == 10'h2ef ? _GEN_3690 : _GEN_3689; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3692 = ~io_inputBit ? 1'h0 : _GEN_3691; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3693 = _GEN_6085 == 10'h2f0 ? _GEN_3692 : _GEN_3691; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3694 = io_inputBit | _GEN_3693; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3695 = _GEN_6085 == 10'h2f0 ? _GEN_3694 : _GEN_3693; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3696 = ~io_inputBit | _GEN_3695; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3697 = _GEN_6085 == 10'h2f1 ? _GEN_3696 : _GEN_3695; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3698 = io_inputBit ? 1'h0 : _GEN_3697; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3699 = _GEN_6085 == 10'h2f1 ? _GEN_3698 : _GEN_3697; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3700 = ~io_inputBit ? 1'h0 : _GEN_3699; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3701 = _GEN_6085 == 10'h2f2 ? _GEN_3700 : _GEN_3699; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3702 = io_inputBit | _GEN_3701; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3703 = _GEN_6085 == 10'h2f2 ? _GEN_3702 : _GEN_3701; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3704 = ~io_inputBit | _GEN_3703; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3705 = _GEN_6085 == 10'h2f3 ? _GEN_3704 : _GEN_3703; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3706 = io_inputBit ? 1'h0 : _GEN_3705; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3707 = _GEN_6085 == 10'h2f3 ? _GEN_3706 : _GEN_3705; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3708 = ~io_inputBit ? 1'h0 : _GEN_3707; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3709 = _GEN_6085 == 10'h2f4 ? _GEN_3708 : _GEN_3707; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3710 = io_inputBit | _GEN_3709; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3711 = _GEN_6085 == 10'h2f4 ? _GEN_3710 : _GEN_3709; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3712 = ~io_inputBit | _GEN_3711; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3713 = _GEN_6085 == 10'h2f5 ? _GEN_3712 : _GEN_3711; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3714 = io_inputBit ? 1'h0 : _GEN_3713; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3715 = _GEN_6085 == 10'h2f5 ? _GEN_3714 : _GEN_3713; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3716 = ~io_inputBit ? 1'h0 : _GEN_3715; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3717 = _GEN_6085 == 10'h2f6 ? _GEN_3716 : _GEN_3715; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3718 = io_inputBit | _GEN_3717; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3719 = _GEN_6085 == 10'h2f6 ? _GEN_3718 : _GEN_3717; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3720 = ~io_inputBit | _GEN_3719; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3721 = _GEN_6085 == 10'h2f7 ? _GEN_3720 : _GEN_3719; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3722 = io_inputBit ? 1'h0 : _GEN_3721; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3723 = _GEN_6085 == 10'h2f7 ? _GEN_3722 : _GEN_3721; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3724 = ~io_inputBit ? 1'h0 : _GEN_3723; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3725 = _GEN_6085 == 10'h2f8 ? _GEN_3724 : _GEN_3723; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3726 = io_inputBit | _GEN_3725; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3727 = _GEN_6085 == 10'h2f8 ? _GEN_3726 : _GEN_3725; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3728 = ~io_inputBit | _GEN_3727; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3729 = _GEN_6085 == 10'h2f9 ? _GEN_3728 : _GEN_3727; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3730 = io_inputBit ? 1'h0 : _GEN_3729; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3731 = _GEN_6085 == 10'h2f9 ? _GEN_3730 : _GEN_3729; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3732 = ~io_inputBit ? 1'h0 : _GEN_3731; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3733 = _GEN_6085 == 10'h2fa ? _GEN_3732 : _GEN_3731; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3734 = io_inputBit | _GEN_3733; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3735 = _GEN_6085 == 10'h2fa ? _GEN_3734 : _GEN_3733; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3736 = ~io_inputBit | _GEN_3735; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3737 = _GEN_6085 == 10'h2fb ? _GEN_3736 : _GEN_3735; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3738 = io_inputBit ? 1'h0 : _GEN_3737; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3739 = _GEN_6085 == 10'h2fb ? _GEN_3738 : _GEN_3737; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3740 = ~io_inputBit ? 1'h0 : _GEN_3739; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3741 = _GEN_6085 == 10'h2fc ? _GEN_3740 : _GEN_3739; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3742 = io_inputBit | _GEN_3741; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3743 = _GEN_6085 == 10'h2fc ? _GEN_3742 : _GEN_3741; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3744 = ~io_inputBit | _GEN_3743; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3745 = _GEN_6085 == 10'h2fd ? _GEN_3744 : _GEN_3743; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3746 = io_inputBit ? 1'h0 : _GEN_3745; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3747 = _GEN_6085 == 10'h2fd ? _GEN_3746 : _GEN_3745; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3748 = ~io_inputBit ? 1'h0 : _GEN_3747; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3749 = _GEN_6085 == 10'h2fe ? _GEN_3748 : _GEN_3747; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3750 = io_inputBit | _GEN_3749; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3751 = _GEN_6085 == 10'h2fe ? _GEN_3750 : _GEN_3749; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3752 = ~io_inputBit | _GEN_3751; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3753 = _GEN_6085 == 10'h2ff ? _GEN_3752 : _GEN_3751; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3754 = io_inputBit ? 1'h0 : _GEN_3753; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3755 = _GEN_6085 == 10'h2ff ? _GEN_3754 : _GEN_3753; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3756 = ~io_inputBit ? 1'h0 : _GEN_3755; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3757 = _GEN_6085 == 10'h300 ? _GEN_3756 : _GEN_3755; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3758 = io_inputBit | _GEN_3757; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3759 = _GEN_6085 == 10'h300 ? _GEN_3758 : _GEN_3757; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3760 = ~io_inputBit | _GEN_3759; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3761 = _GEN_6085 == 10'h301 ? _GEN_3760 : _GEN_3759; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3762 = io_inputBit ? 1'h0 : _GEN_3761; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3763 = _GEN_6085 == 10'h301 ? _GEN_3762 : _GEN_3761; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3764 = ~io_inputBit ? 1'h0 : _GEN_3763; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3765 = _GEN_6085 == 10'h302 ? _GEN_3764 : _GEN_3763; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3766 = io_inputBit | _GEN_3765; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3767 = _GEN_6085 == 10'h302 ? _GEN_3766 : _GEN_3765; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3768 = ~io_inputBit | _GEN_3767; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3769 = _GEN_6085 == 10'h303 ? _GEN_3768 : _GEN_3767; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3770 = io_inputBit ? 1'h0 : _GEN_3769; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3771 = _GEN_6085 == 10'h303 ? _GEN_3770 : _GEN_3769; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3772 = ~io_inputBit ? 1'h0 : _GEN_3771; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3773 = _GEN_6085 == 10'h304 ? _GEN_3772 : _GEN_3771; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3774 = io_inputBit | _GEN_3773; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3775 = _GEN_6085 == 10'h304 ? _GEN_3774 : _GEN_3773; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3776 = ~io_inputBit | _GEN_3775; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3777 = _GEN_6085 == 10'h305 ? _GEN_3776 : _GEN_3775; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3778 = io_inputBit ? 1'h0 : _GEN_3777; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3779 = _GEN_6085 == 10'h305 ? _GEN_3778 : _GEN_3777; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3780 = ~io_inputBit ? 1'h0 : _GEN_3779; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3781 = _GEN_6085 == 10'h306 ? _GEN_3780 : _GEN_3779; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3782 = io_inputBit | _GEN_3781; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3783 = _GEN_6085 == 10'h306 ? _GEN_3782 : _GEN_3781; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3784 = ~io_inputBit | _GEN_3783; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3785 = _GEN_6085 == 10'h307 ? _GEN_3784 : _GEN_3783; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3786 = io_inputBit ? 1'h0 : _GEN_3785; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3787 = _GEN_6085 == 10'h307 ? _GEN_3786 : _GEN_3785; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3788 = ~io_inputBit ? 1'h0 : _GEN_3787; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3789 = _GEN_6085 == 10'h308 ? _GEN_3788 : _GEN_3787; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3790 = io_inputBit | _GEN_3789; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3791 = _GEN_6085 == 10'h308 ? _GEN_3790 : _GEN_3789; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3792 = ~io_inputBit | _GEN_3791; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3793 = _GEN_6085 == 10'h309 ? _GEN_3792 : _GEN_3791; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3794 = io_inputBit ? 1'h0 : _GEN_3793; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3795 = _GEN_6085 == 10'h309 ? _GEN_3794 : _GEN_3793; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3796 = ~io_inputBit ? 1'h0 : _GEN_3795; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3797 = _GEN_6085 == 10'h30a ? _GEN_3796 : _GEN_3795; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3798 = io_inputBit | _GEN_3797; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3799 = _GEN_6085 == 10'h30a ? _GEN_3798 : _GEN_3797; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3800 = ~io_inputBit | _GEN_3799; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3801 = _GEN_6085 == 10'h30b ? _GEN_3800 : _GEN_3799; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3802 = io_inputBit ? 1'h0 : _GEN_3801; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3803 = _GEN_6085 == 10'h30b ? _GEN_3802 : _GEN_3801; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3804 = ~io_inputBit ? 1'h0 : _GEN_3803; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3805 = _GEN_6085 == 10'h30c ? _GEN_3804 : _GEN_3803; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3806 = io_inputBit | _GEN_3805; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3807 = _GEN_6085 == 10'h30c ? _GEN_3806 : _GEN_3805; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3808 = ~io_inputBit | _GEN_3807; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3809 = _GEN_6085 == 10'h30d ? _GEN_3808 : _GEN_3807; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3810 = io_inputBit ? 1'h0 : _GEN_3809; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3811 = _GEN_6085 == 10'h30d ? _GEN_3810 : _GEN_3809; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3812 = ~io_inputBit ? 1'h0 : _GEN_3811; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3813 = _GEN_6085 == 10'h30e ? _GEN_3812 : _GEN_3811; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3814 = io_inputBit | _GEN_3813; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3815 = _GEN_6085 == 10'h30e ? _GEN_3814 : _GEN_3813; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3816 = ~io_inputBit | _GEN_3815; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3817 = _GEN_6085 == 10'h30f ? _GEN_3816 : _GEN_3815; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3818 = io_inputBit ? 1'h0 : _GEN_3817; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3819 = _GEN_6085 == 10'h30f ? _GEN_3818 : _GEN_3817; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3820 = ~io_inputBit ? 1'h0 : _GEN_3819; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3821 = _GEN_6085 == 10'h310 ? _GEN_3820 : _GEN_3819; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3822 = io_inputBit | _GEN_3821; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3823 = _GEN_6085 == 10'h310 ? _GEN_3822 : _GEN_3821; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3824 = ~io_inputBit | _GEN_3823; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3825 = _GEN_6085 == 10'h311 ? _GEN_3824 : _GEN_3823; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3826 = io_inputBit ? 1'h0 : _GEN_3825; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3827 = _GEN_6085 == 10'h311 ? _GEN_3826 : _GEN_3825; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3828 = ~io_inputBit ? 1'h0 : _GEN_2831; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3829 = i == 8'h1 ? _GEN_3828 : _GEN_2831; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3830 = io_inputBit ? 1'h0 : _GEN_3829; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3831 = i == 8'h2 ? _GEN_3830 : _GEN_3829; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3832 = io_inputBit ? 1'h0 : _GEN_3831; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3833 = i == 8'h5 ? _GEN_3832 : _GEN_3831; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3834 = ~io_inputBit ? 1'h0 : _GEN_3833; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3835 = i == 8'h9 ? _GEN_3834 : _GEN_3833; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3836 = io_inputBit ? 1'h0 : _GEN_3835; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3837 = i == 8'hb ? _GEN_3836 : _GEN_3835; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3838 = ~io_inputBit ? 1'h0 : _GEN_3837; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3839 = i == 8'h29 ? _GEN_3838 : _GEN_3837; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3840 = io_inputBit ? 1'h0 : _GEN_3839; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3841 = i == 8'h30 ? _GEN_3840 : _GEN_3839; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3842 = ~io_inputBit ? 1'h0 : _GEN_3841; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3843 = i == 8'h54 ? _GEN_3842 : _GEN_3841; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3844 = io_inputBit ? 1'h0 : _GEN_3843; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3845 = i == 8'h61 ? _GEN_3844 : _GEN_3843; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3846 = ~io_inputBit ? 1'h0 : _GEN_3845; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3847 = i == 8'haa ? _GEN_3846 : _GEN_3845; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3848 = ~io_inputBit ? 1'h0 : _GEN_3847; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3849 = _GEN_6084 == 9'h156 ? _GEN_3848 : _GEN_3847; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3850 = io_inputBit ? 1'h0 : _GEN_3849; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3851 = _GEN_6084 == 9'h188 ? _GEN_3850 : _GEN_3849; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3852 = ~io_inputBit ? 1'h0 : _GEN_3851; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3853 = _GEN_6085 == 10'h2ae ? _GEN_3852 : _GEN_3851; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3854 = io_inputBit | _GEN_3853; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3855 = _GEN_6085 == 10'h2ae ? _GEN_3854 : _GEN_3853; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3856 = ~io_inputBit ? 1'h0 : _GEN_3855; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3857 = _GEN_6085 == 10'h2af ? _GEN_3856 : _GEN_3855; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3858 = io_inputBit | _GEN_3857; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3859 = _GEN_6085 == 10'h2af ? _GEN_3858 : _GEN_3857; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3860 = ~io_inputBit ? 1'h0 : _GEN_3859; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3861 = _GEN_6085 == 10'h2b0 ? _GEN_3860 : _GEN_3859; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3862 = io_inputBit | _GEN_3861; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3863 = _GEN_6085 == 10'h2b0 ? _GEN_3862 : _GEN_3861; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3864 = ~io_inputBit ? 1'h0 : _GEN_3863; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3865 = _GEN_6085 == 10'h2b1 ? _GEN_3864 : _GEN_3863; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3866 = io_inputBit | _GEN_3865; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3867 = _GEN_6085 == 10'h2b1 ? _GEN_3866 : _GEN_3865; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3868 = ~io_inputBit ? 1'h0 : _GEN_3867; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3869 = _GEN_6085 == 10'h2b2 ? _GEN_3868 : _GEN_3867; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3870 = io_inputBit | _GEN_3869; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3871 = _GEN_6085 == 10'h2b2 ? _GEN_3870 : _GEN_3869; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3872 = ~io_inputBit ? 1'h0 : _GEN_3871; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3873 = _GEN_6085 == 10'h2b3 ? _GEN_3872 : _GEN_3871; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3874 = io_inputBit | _GEN_3873; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3875 = _GEN_6085 == 10'h2b3 ? _GEN_3874 : _GEN_3873; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3876 = ~io_inputBit ? 1'h0 : _GEN_3875; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3877 = _GEN_6085 == 10'h2b4 ? _GEN_3876 : _GEN_3875; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3878 = io_inputBit | _GEN_3877; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3879 = _GEN_6085 == 10'h2b4 ? _GEN_3878 : _GEN_3877; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3880 = ~io_inputBit ? 1'h0 : _GEN_3879; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3881 = _GEN_6085 == 10'h2b5 ? _GEN_3880 : _GEN_3879; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3882 = io_inputBit | _GEN_3881; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3883 = _GEN_6085 == 10'h2b5 ? _GEN_3882 : _GEN_3881; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3884 = ~io_inputBit ? 1'h0 : _GEN_3883; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3885 = _GEN_6085 == 10'h2b6 ? _GEN_3884 : _GEN_3883; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3886 = io_inputBit | _GEN_3885; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3887 = _GEN_6085 == 10'h2b6 ? _GEN_3886 : _GEN_3885; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3888 = ~io_inputBit ? 1'h0 : _GEN_3887; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3889 = _GEN_6085 == 10'h2b7 ? _GEN_3888 : _GEN_3887; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3890 = io_inputBit | _GEN_3889; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3891 = _GEN_6085 == 10'h2b7 ? _GEN_3890 : _GEN_3889; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3892 = ~io_inputBit ? 1'h0 : _GEN_3891; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3893 = _GEN_6085 == 10'h2b8 ? _GEN_3892 : _GEN_3891; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3894 = io_inputBit | _GEN_3893; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3895 = _GEN_6085 == 10'h2b8 ? _GEN_3894 : _GEN_3893; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3896 = ~io_inputBit ? 1'h0 : _GEN_3895; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3897 = _GEN_6085 == 10'h2b9 ? _GEN_3896 : _GEN_3895; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3898 = io_inputBit | _GEN_3897; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3899 = _GEN_6085 == 10'h2b9 ? _GEN_3898 : _GEN_3897; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3900 = ~io_inputBit ? 1'h0 : _GEN_3899; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3901 = _GEN_6085 == 10'h2ba ? _GEN_3900 : _GEN_3899; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3902 = io_inputBit | _GEN_3901; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3903 = _GEN_6085 == 10'h2ba ? _GEN_3902 : _GEN_3901; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3904 = ~io_inputBit ? 1'h0 : _GEN_3903; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3905 = _GEN_6085 == 10'h2bb ? _GEN_3904 : _GEN_3903; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3906 = io_inputBit | _GEN_3905; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3907 = _GEN_6085 == 10'h2bb ? _GEN_3906 : _GEN_3905; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3908 = ~io_inputBit ? 1'h0 : _GEN_3907; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3909 = _GEN_6085 == 10'h2bc ? _GEN_3908 : _GEN_3907; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3910 = io_inputBit | _GEN_3909; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3911 = _GEN_6085 == 10'h2bc ? _GEN_3910 : _GEN_3909; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3912 = ~io_inputBit ? 1'h0 : _GEN_3911; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3913 = _GEN_6085 == 10'h2bd ? _GEN_3912 : _GEN_3911; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3914 = io_inputBit | _GEN_3913; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3915 = _GEN_6085 == 10'h2bd ? _GEN_3914 : _GEN_3913; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3916 = ~io_inputBit ? 1'h0 : _GEN_3915; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3917 = _GEN_6085 == 10'h2be ? _GEN_3916 : _GEN_3915; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3918 = io_inputBit | _GEN_3917; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3919 = _GEN_6085 == 10'h2be ? _GEN_3918 : _GEN_3917; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3920 = ~io_inputBit ? 1'h0 : _GEN_3919; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3921 = _GEN_6085 == 10'h2bf ? _GEN_3920 : _GEN_3919; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3922 = io_inputBit | _GEN_3921; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3923 = _GEN_6085 == 10'h2bf ? _GEN_3922 : _GEN_3921; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3924 = ~io_inputBit ? 1'h0 : _GEN_3923; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3925 = _GEN_6085 == 10'h2c0 ? _GEN_3924 : _GEN_3923; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3926 = io_inputBit | _GEN_3925; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3927 = _GEN_6085 == 10'h2c0 ? _GEN_3926 : _GEN_3925; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3928 = ~io_inputBit ? 1'h0 : _GEN_3927; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3929 = _GEN_6085 == 10'h2c1 ? _GEN_3928 : _GEN_3927; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3930 = io_inputBit | _GEN_3929; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3931 = _GEN_6085 == 10'h2c1 ? _GEN_3930 : _GEN_3929; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3932 = ~io_inputBit ? 1'h0 : _GEN_3931; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3933 = _GEN_6085 == 10'h2c2 ? _GEN_3932 : _GEN_3931; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3934 = io_inputBit | _GEN_3933; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3935 = _GEN_6085 == 10'h2c2 ? _GEN_3934 : _GEN_3933; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3936 = ~io_inputBit ? 1'h0 : _GEN_3935; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3937 = _GEN_6085 == 10'h2c3 ? _GEN_3936 : _GEN_3935; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3938 = io_inputBit | _GEN_3937; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3939 = _GEN_6085 == 10'h2c3 ? _GEN_3938 : _GEN_3937; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3940 = ~io_inputBit ? 1'h0 : _GEN_3939; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3941 = _GEN_6085 == 10'h2c4 ? _GEN_3940 : _GEN_3939; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3942 = io_inputBit | _GEN_3941; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3943 = _GEN_6085 == 10'h2c4 ? _GEN_3942 : _GEN_3941; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3944 = ~io_inputBit ? 1'h0 : _GEN_3943; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3945 = _GEN_6085 == 10'h2c5 ? _GEN_3944 : _GEN_3943; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3946 = io_inputBit | _GEN_3945; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3947 = _GEN_6085 == 10'h2c5 ? _GEN_3946 : _GEN_3945; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3948 = ~io_inputBit ? 1'h0 : _GEN_3947; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3949 = _GEN_6085 == 10'h2c6 ? _GEN_3948 : _GEN_3947; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3950 = io_inputBit | _GEN_3949; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3951 = _GEN_6085 == 10'h2c6 ? _GEN_3950 : _GEN_3949; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3952 = ~io_inputBit ? 1'h0 : _GEN_3951; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3953 = _GEN_6085 == 10'h2c7 ? _GEN_3952 : _GEN_3951; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3954 = io_inputBit | _GEN_3953; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3955 = _GEN_6085 == 10'h2c7 ? _GEN_3954 : _GEN_3953; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3956 = ~io_inputBit ? 1'h0 : _GEN_3955; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3957 = _GEN_6085 == 10'h2c8 ? _GEN_3956 : _GEN_3955; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3958 = io_inputBit | _GEN_3957; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3959 = _GEN_6085 == 10'h2c8 ? _GEN_3958 : _GEN_3957; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3960 = ~io_inputBit ? 1'h0 : _GEN_3959; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3961 = _GEN_6085 == 10'h2c9 ? _GEN_3960 : _GEN_3959; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3962 = io_inputBit | _GEN_3961; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3963 = _GEN_6085 == 10'h2c9 ? _GEN_3962 : _GEN_3961; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3964 = ~io_inputBit ? 1'h0 : _GEN_3963; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3965 = _GEN_6085 == 10'h2ca ? _GEN_3964 : _GEN_3963; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3966 = io_inputBit | _GEN_3965; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3967 = _GEN_6085 == 10'h2ca ? _GEN_3966 : _GEN_3965; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3968 = ~io_inputBit ? 1'h0 : _GEN_3967; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3969 = _GEN_6085 == 10'h2cb ? _GEN_3968 : _GEN_3967; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3970 = io_inputBit | _GEN_3969; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3971 = _GEN_6085 == 10'h2cb ? _GEN_3970 : _GEN_3969; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3972 = ~io_inputBit ? 1'h0 : _GEN_3971; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3973 = _GEN_6085 == 10'h2cc ? _GEN_3972 : _GEN_3971; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3974 = io_inputBit | _GEN_3973; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3975 = _GEN_6085 == 10'h2cc ? _GEN_3974 : _GEN_3973; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3976 = ~io_inputBit ? 1'h0 : _GEN_3975; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3977 = _GEN_6085 == 10'h2cd ? _GEN_3976 : _GEN_3975; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3978 = io_inputBit | _GEN_3977; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3979 = _GEN_6085 == 10'h2cd ? _GEN_3978 : _GEN_3977; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3980 = ~io_inputBit ? 1'h0 : _GEN_3979; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3981 = _GEN_6085 == 10'h2ce ? _GEN_3980 : _GEN_3979; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3982 = io_inputBit | _GEN_3981; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3983 = _GEN_6085 == 10'h2ce ? _GEN_3982 : _GEN_3981; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3984 = ~io_inputBit ? 1'h0 : _GEN_3983; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3985 = _GEN_6085 == 10'h2cf ? _GEN_3984 : _GEN_3983; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3986 = io_inputBit | _GEN_3985; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3987 = _GEN_6085 == 10'h2cf ? _GEN_3986 : _GEN_3985; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3988 = ~io_inputBit ? 1'h0 : _GEN_3987; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3989 = _GEN_6085 == 10'h2d0 ? _GEN_3988 : _GEN_3987; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3990 = io_inputBit | _GEN_3989; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3991 = _GEN_6085 == 10'h2d0 ? _GEN_3990 : _GEN_3989; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3992 = ~io_inputBit ? 1'h0 : _GEN_3991; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3993 = _GEN_6085 == 10'h2d1 ? _GEN_3992 : _GEN_3991; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3994 = io_inputBit | _GEN_3993; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3995 = _GEN_6085 == 10'h2d1 ? _GEN_3994 : _GEN_3993; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3996 = ~io_inputBit ? 1'h0 : _GEN_3995; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3997 = _GEN_6085 == 10'h2d2 ? _GEN_3996 : _GEN_3995; // @[lut_mem_online.scala 235:34]
  wire  _GEN_3998 = io_inputBit | _GEN_3997; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_3999 = _GEN_6085 == 10'h2d2 ? _GEN_3998 : _GEN_3997; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4000 = ~io_inputBit ? 1'h0 : _GEN_3999; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4001 = _GEN_6085 == 10'h2d3 ? _GEN_4000 : _GEN_3999; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4002 = io_inputBit | _GEN_4001; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4003 = _GEN_6085 == 10'h2d3 ? _GEN_4002 : _GEN_4001; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4004 = ~io_inputBit ? 1'h0 : _GEN_4003; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4005 = _GEN_6085 == 10'h2d4 ? _GEN_4004 : _GEN_4003; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4006 = io_inputBit | _GEN_4005; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4007 = _GEN_6085 == 10'h2d4 ? _GEN_4006 : _GEN_4005; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4008 = ~io_inputBit ? 1'h0 : _GEN_4007; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4009 = _GEN_6085 == 10'h2d5 ? _GEN_4008 : _GEN_4007; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4010 = io_inputBit | _GEN_4009; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4011 = _GEN_6085 == 10'h2d5 ? _GEN_4010 : _GEN_4009; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4012 = ~io_inputBit ? 1'h0 : _GEN_4011; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4013 = _GEN_6085 == 10'h2d6 ? _GEN_4012 : _GEN_4011; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4014 = io_inputBit | _GEN_4013; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4015 = _GEN_6085 == 10'h2d6 ? _GEN_4014 : _GEN_4013; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4016 = ~io_inputBit ? 1'h0 : _GEN_4015; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4017 = _GEN_6085 == 10'h2d7 ? _GEN_4016 : _GEN_4015; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4018 = io_inputBit | _GEN_4017; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4019 = _GEN_6085 == 10'h2d7 ? _GEN_4018 : _GEN_4017; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4020 = ~io_inputBit ? 1'h0 : _GEN_4019; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4021 = _GEN_6085 == 10'h2d8 ? _GEN_4020 : _GEN_4019; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4022 = io_inputBit | _GEN_4021; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4023 = _GEN_6085 == 10'h2d8 ? _GEN_4022 : _GEN_4021; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4024 = ~io_inputBit ? 1'h0 : _GEN_4023; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4025 = _GEN_6085 == 10'h2d9 ? _GEN_4024 : _GEN_4023; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4026 = io_inputBit | _GEN_4025; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4027 = _GEN_6085 == 10'h2d9 ? _GEN_4026 : _GEN_4025; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4028 = ~io_inputBit ? 1'h0 : _GEN_4027; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4029 = _GEN_6085 == 10'h2da ? _GEN_4028 : _GEN_4027; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4030 = io_inputBit | _GEN_4029; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4031 = _GEN_6085 == 10'h2da ? _GEN_4030 : _GEN_4029; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4032 = ~io_inputBit ? 1'h0 : _GEN_4031; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4033 = _GEN_6085 == 10'h2db ? _GEN_4032 : _GEN_4031; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4034 = io_inputBit | _GEN_4033; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4035 = _GEN_6085 == 10'h2db ? _GEN_4034 : _GEN_4033; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4036 = ~io_inputBit ? 1'h0 : _GEN_4035; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4037 = _GEN_6085 == 10'h2dc ? _GEN_4036 : _GEN_4035; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4038 = io_inputBit | _GEN_4037; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4039 = _GEN_6085 == 10'h2dc ? _GEN_4038 : _GEN_4037; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4040 = ~io_inputBit ? 1'h0 : _GEN_4039; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4041 = _GEN_6085 == 10'h2dd ? _GEN_4040 : _GEN_4039; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4042 = io_inputBit | _GEN_4041; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4043 = _GEN_6085 == 10'h2dd ? _GEN_4042 : _GEN_4041; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4044 = ~io_inputBit ? 1'h0 : _GEN_4043; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4045 = _GEN_6085 == 10'h2de ? _GEN_4044 : _GEN_4043; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4046 = io_inputBit | _GEN_4045; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4047 = _GEN_6085 == 10'h2de ? _GEN_4046 : _GEN_4045; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4048 = ~io_inputBit ? 1'h0 : _GEN_4047; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4049 = _GEN_6085 == 10'h2df ? _GEN_4048 : _GEN_4047; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4050 = io_inputBit | _GEN_4049; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4051 = _GEN_6085 == 10'h2df ? _GEN_4050 : _GEN_4049; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4052 = ~io_inputBit ? 1'h0 : _GEN_4051; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4053 = _GEN_6085 == 10'h2e0 ? _GEN_4052 : _GEN_4051; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4054 = io_inputBit | _GEN_4053; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4055 = _GEN_6085 == 10'h2e0 ? _GEN_4054 : _GEN_4053; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4056 = ~io_inputBit ? 1'h0 : _GEN_4055; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4057 = _GEN_6085 == 10'h2e1 ? _GEN_4056 : _GEN_4055; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4058 = io_inputBit | _GEN_4057; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4059 = _GEN_6085 == 10'h2e1 ? _GEN_4058 : _GEN_4057; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4060 = ~io_inputBit ? 1'h0 : _GEN_4059; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4061 = _GEN_6085 == 10'h2e2 ? _GEN_4060 : _GEN_4059; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4062 = io_inputBit | _GEN_4061; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4063 = _GEN_6085 == 10'h2e2 ? _GEN_4062 : _GEN_4061; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4064 = ~io_inputBit ? 1'h0 : _GEN_4063; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4065 = _GEN_6085 == 10'h2e3 ? _GEN_4064 : _GEN_4063; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4066 = io_inputBit | _GEN_4065; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4067 = _GEN_6085 == 10'h2e3 ? _GEN_4066 : _GEN_4065; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4068 = ~io_inputBit ? 1'h0 : _GEN_4067; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4069 = _GEN_6085 == 10'h2e4 ? _GEN_4068 : _GEN_4067; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4070 = io_inputBit | _GEN_4069; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4071 = _GEN_6085 == 10'h2e4 ? _GEN_4070 : _GEN_4069; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4072 = ~io_inputBit ? 1'h0 : _GEN_4071; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4073 = _GEN_6085 == 10'h2e5 ? _GEN_4072 : _GEN_4071; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4074 = io_inputBit | _GEN_4073; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4075 = _GEN_6085 == 10'h2e5 ? _GEN_4074 : _GEN_4073; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4076 = ~io_inputBit ? 1'h0 : _GEN_4075; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4077 = _GEN_6085 == 10'h2e6 ? _GEN_4076 : _GEN_4075; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4078 = io_inputBit | _GEN_4077; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4079 = _GEN_6085 == 10'h2e6 ? _GEN_4078 : _GEN_4077; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4080 = ~io_inputBit ? 1'h0 : _GEN_4079; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4081 = _GEN_6085 == 10'h2e7 ? _GEN_4080 : _GEN_4079; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4082 = io_inputBit | _GEN_4081; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4083 = _GEN_6085 == 10'h2e7 ? _GEN_4082 : _GEN_4081; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4084 = ~io_inputBit ? 1'h0 : _GEN_4083; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4085 = _GEN_6085 == 10'h2e8 ? _GEN_4084 : _GEN_4083; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4086 = io_inputBit | _GEN_4085; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4087 = _GEN_6085 == 10'h2e8 ? _GEN_4086 : _GEN_4085; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4088 = ~io_inputBit ? 1'h0 : _GEN_4087; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4089 = _GEN_6085 == 10'h2e9 ? _GEN_4088 : _GEN_4087; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4090 = io_inputBit | _GEN_4089; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4091 = _GEN_6085 == 10'h2e9 ? _GEN_4090 : _GEN_4089; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4092 = ~io_inputBit ? 1'h0 : _GEN_4091; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4093 = _GEN_6085 == 10'h2ea ? _GEN_4092 : _GEN_4091; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4094 = io_inputBit | _GEN_4093; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4095 = _GEN_6085 == 10'h2ea ? _GEN_4094 : _GEN_4093; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4096 = ~io_inputBit ? 1'h0 : _GEN_4095; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4097 = _GEN_6085 == 10'h2eb ? _GEN_4096 : _GEN_4095; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4098 = io_inputBit | _GEN_4097; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4099 = _GEN_6085 == 10'h2eb ? _GEN_4098 : _GEN_4097; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4100 = ~io_inputBit ? 1'h0 : _GEN_4099; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4101 = _GEN_6085 == 10'h2ec ? _GEN_4100 : _GEN_4099; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4102 = io_inputBit | _GEN_4101; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4103 = _GEN_6085 == 10'h2ec ? _GEN_4102 : _GEN_4101; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4104 = ~io_inputBit ? 1'h0 : _GEN_4103; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4105 = _GEN_6085 == 10'h2ed ? _GEN_4104 : _GEN_4103; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4106 = io_inputBit | _GEN_4105; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4107 = _GEN_6085 == 10'h2ed ? _GEN_4106 : _GEN_4105; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4108 = ~io_inputBit ? 1'h0 : _GEN_4107; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4109 = _GEN_6085 == 10'h2ee ? _GEN_4108 : _GEN_4107; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4110 = io_inputBit | _GEN_4109; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4111 = _GEN_6085 == 10'h2ee ? _GEN_4110 : _GEN_4109; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4112 = ~io_inputBit ? 1'h0 : _GEN_4111; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4113 = _GEN_6085 == 10'h2ef ? _GEN_4112 : _GEN_4111; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4114 = io_inputBit | _GEN_4113; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4115 = _GEN_6085 == 10'h2ef ? _GEN_4114 : _GEN_4113; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4116 = ~io_inputBit ? 1'h0 : _GEN_4115; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4117 = _GEN_6085 == 10'h2f0 ? _GEN_4116 : _GEN_4115; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4118 = io_inputBit | _GEN_4117; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4119 = _GEN_6085 == 10'h2f0 ? _GEN_4118 : _GEN_4117; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4120 = ~io_inputBit ? 1'h0 : _GEN_4119; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4121 = _GEN_6085 == 10'h2f1 ? _GEN_4120 : _GEN_4119; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4122 = io_inputBit | _GEN_4121; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4123 = _GEN_6085 == 10'h2f1 ? _GEN_4122 : _GEN_4121; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4124 = ~io_inputBit ? 1'h0 : _GEN_4123; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4125 = _GEN_6085 == 10'h2f2 ? _GEN_4124 : _GEN_4123; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4126 = io_inputBit | _GEN_4125; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4127 = _GEN_6085 == 10'h2f2 ? _GEN_4126 : _GEN_4125; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4128 = ~io_inputBit ? 1'h0 : _GEN_4127; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4129 = _GEN_6085 == 10'h2f3 ? _GEN_4128 : _GEN_4127; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4130 = io_inputBit | _GEN_4129; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4131 = _GEN_6085 == 10'h2f3 ? _GEN_4130 : _GEN_4129; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4132 = ~io_inputBit ? 1'h0 : _GEN_4131; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4133 = _GEN_6085 == 10'h2f4 ? _GEN_4132 : _GEN_4131; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4134 = io_inputBit | _GEN_4133; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4135 = _GEN_6085 == 10'h2f4 ? _GEN_4134 : _GEN_4133; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4136 = ~io_inputBit ? 1'h0 : _GEN_4135; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4137 = _GEN_6085 == 10'h2f5 ? _GEN_4136 : _GEN_4135; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4138 = io_inputBit | _GEN_4137; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4139 = _GEN_6085 == 10'h2f5 ? _GEN_4138 : _GEN_4137; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4140 = ~io_inputBit ? 1'h0 : _GEN_4139; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4141 = _GEN_6085 == 10'h2f6 ? _GEN_4140 : _GEN_4139; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4142 = io_inputBit | _GEN_4141; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4143 = _GEN_6085 == 10'h2f6 ? _GEN_4142 : _GEN_4141; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4144 = ~io_inputBit ? 1'h0 : _GEN_4143; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4145 = _GEN_6085 == 10'h2f7 ? _GEN_4144 : _GEN_4143; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4146 = io_inputBit | _GEN_4145; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4147 = _GEN_6085 == 10'h2f7 ? _GEN_4146 : _GEN_4145; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4148 = ~io_inputBit ? 1'h0 : _GEN_4147; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4149 = _GEN_6085 == 10'h2f8 ? _GEN_4148 : _GEN_4147; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4150 = io_inputBit | _GEN_4149; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4151 = _GEN_6085 == 10'h2f8 ? _GEN_4150 : _GEN_4149; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4152 = ~io_inputBit ? 1'h0 : _GEN_4151; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4153 = _GEN_6085 == 10'h2f9 ? _GEN_4152 : _GEN_4151; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4154 = io_inputBit | _GEN_4153; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4155 = _GEN_6085 == 10'h2f9 ? _GEN_4154 : _GEN_4153; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4156 = ~io_inputBit ? 1'h0 : _GEN_4155; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4157 = _GEN_6085 == 10'h2fa ? _GEN_4156 : _GEN_4155; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4158 = io_inputBit | _GEN_4157; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4159 = _GEN_6085 == 10'h2fa ? _GEN_4158 : _GEN_4157; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4160 = ~io_inputBit ? 1'h0 : _GEN_4159; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4161 = _GEN_6085 == 10'h2fb ? _GEN_4160 : _GEN_4159; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4162 = io_inputBit | _GEN_4161; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4163 = _GEN_6085 == 10'h2fb ? _GEN_4162 : _GEN_4161; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4164 = ~io_inputBit ? 1'h0 : _GEN_4163; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4165 = _GEN_6085 == 10'h2fc ? _GEN_4164 : _GEN_4163; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4166 = io_inputBit | _GEN_4165; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4167 = _GEN_6085 == 10'h2fc ? _GEN_4166 : _GEN_4165; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4168 = ~io_inputBit ? 1'h0 : _GEN_4167; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4169 = _GEN_6085 == 10'h2fd ? _GEN_4168 : _GEN_4167; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4170 = io_inputBit | _GEN_4169; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4171 = _GEN_6085 == 10'h2fd ? _GEN_4170 : _GEN_4169; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4172 = ~io_inputBit ? 1'h0 : _GEN_4171; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4173 = _GEN_6085 == 10'h2fe ? _GEN_4172 : _GEN_4171; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4174 = io_inputBit | _GEN_4173; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4175 = _GEN_6085 == 10'h2fe ? _GEN_4174 : _GEN_4173; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4176 = ~io_inputBit ? 1'h0 : _GEN_4175; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4177 = _GEN_6085 == 10'h2ff ? _GEN_4176 : _GEN_4175; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4178 = io_inputBit | _GEN_4177; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4179 = _GEN_6085 == 10'h2ff ? _GEN_4178 : _GEN_4177; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4180 = ~io_inputBit ? 1'h0 : _GEN_4179; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4181 = _GEN_6085 == 10'h300 ? _GEN_4180 : _GEN_4179; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4182 = io_inputBit | _GEN_4181; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4183 = _GEN_6085 == 10'h300 ? _GEN_4182 : _GEN_4181; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4184 = ~io_inputBit ? 1'h0 : _GEN_4183; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4185 = _GEN_6085 == 10'h301 ? _GEN_4184 : _GEN_4183; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4186 = io_inputBit | _GEN_4185; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4187 = _GEN_6085 == 10'h301 ? _GEN_4186 : _GEN_4185; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4188 = ~io_inputBit ? 1'h0 : _GEN_4187; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4189 = _GEN_6085 == 10'h302 ? _GEN_4188 : _GEN_4187; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4190 = io_inputBit | _GEN_4189; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4191 = _GEN_6085 == 10'h302 ? _GEN_4190 : _GEN_4189; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4192 = ~io_inputBit ? 1'h0 : _GEN_4191; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4193 = _GEN_6085 == 10'h303 ? _GEN_4192 : _GEN_4191; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4194 = io_inputBit | _GEN_4193; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4195 = _GEN_6085 == 10'h303 ? _GEN_4194 : _GEN_4193; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4196 = ~io_inputBit ? 1'h0 : _GEN_4195; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4197 = _GEN_6085 == 10'h304 ? _GEN_4196 : _GEN_4195; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4198 = io_inputBit | _GEN_4197; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4199 = _GEN_6085 == 10'h304 ? _GEN_4198 : _GEN_4197; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4200 = ~io_inputBit ? 1'h0 : _GEN_4199; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4201 = _GEN_6085 == 10'h305 ? _GEN_4200 : _GEN_4199; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4202 = io_inputBit | _GEN_4201; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4203 = _GEN_6085 == 10'h305 ? _GEN_4202 : _GEN_4201; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4204 = ~io_inputBit ? 1'h0 : _GEN_4203; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4205 = _GEN_6085 == 10'h306 ? _GEN_4204 : _GEN_4203; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4206 = io_inputBit | _GEN_4205; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4207 = _GEN_6085 == 10'h306 ? _GEN_4206 : _GEN_4205; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4208 = ~io_inputBit ? 1'h0 : _GEN_4207; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4209 = _GEN_6085 == 10'h307 ? _GEN_4208 : _GEN_4207; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4210 = io_inputBit | _GEN_4209; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4211 = _GEN_6085 == 10'h307 ? _GEN_4210 : _GEN_4209; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4212 = ~io_inputBit ? 1'h0 : _GEN_4211; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4213 = _GEN_6085 == 10'h308 ? _GEN_4212 : _GEN_4211; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4214 = io_inputBit | _GEN_4213; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4215 = _GEN_6085 == 10'h308 ? _GEN_4214 : _GEN_4213; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4216 = ~io_inputBit ? 1'h0 : _GEN_4215; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4217 = _GEN_6085 == 10'h309 ? _GEN_4216 : _GEN_4215; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4218 = io_inputBit | _GEN_4217; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4219 = _GEN_6085 == 10'h309 ? _GEN_4218 : _GEN_4217; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4220 = ~io_inputBit ? 1'h0 : _GEN_4219; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4221 = _GEN_6085 == 10'h30a ? _GEN_4220 : _GEN_4219; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4222 = io_inputBit | _GEN_4221; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4223 = _GEN_6085 == 10'h30a ? _GEN_4222 : _GEN_4221; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4224 = ~io_inputBit ? 1'h0 : _GEN_4223; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4225 = _GEN_6085 == 10'h30b ? _GEN_4224 : _GEN_4223; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4226 = io_inputBit | _GEN_4225; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4227 = _GEN_6085 == 10'h30b ? _GEN_4226 : _GEN_4225; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4228 = ~io_inputBit ? 1'h0 : _GEN_4227; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4229 = _GEN_6085 == 10'h30c ? _GEN_4228 : _GEN_4227; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4230 = io_inputBit | _GEN_4229; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4231 = _GEN_6085 == 10'h30c ? _GEN_4230 : _GEN_4229; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4232 = ~io_inputBit ? 1'h0 : _GEN_4231; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4233 = _GEN_6085 == 10'h30d ? _GEN_4232 : _GEN_4231; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4234 = io_inputBit | _GEN_4233; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4235 = _GEN_6085 == 10'h30d ? _GEN_4234 : _GEN_4233; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4236 = ~io_inputBit ? 1'h0 : _GEN_4235; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4237 = _GEN_6085 == 10'h30e ? _GEN_4236 : _GEN_4235; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4238 = io_inputBit | _GEN_4237; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4239 = _GEN_6085 == 10'h30e ? _GEN_4238 : _GEN_4237; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4240 = ~io_inputBit ? 1'h0 : _GEN_4239; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4241 = _GEN_6085 == 10'h30f ? _GEN_4240 : _GEN_4239; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4242 = io_inputBit | _GEN_4241; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4243 = _GEN_6085 == 10'h30f ? _GEN_4242 : _GEN_4241; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4244 = ~io_inputBit ? 1'h0 : _GEN_4243; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4245 = _GEN_6085 == 10'h310 ? _GEN_4244 : _GEN_4243; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4246 = io_inputBit | _GEN_4245; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4247 = _GEN_6085 == 10'h310 ? _GEN_4246 : _GEN_4245; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4248 = ~io_inputBit ? 1'h0 : _GEN_4247; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4249 = _GEN_6085 == 10'h311 ? _GEN_4248 : _GEN_4247; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4250 = io_inputBit | _GEN_4249; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4251 = _GEN_6085 == 10'h311 ? _GEN_4250 : _GEN_4249; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4252 = ~io_inputBit ? 1'h0 : _GEN_2863; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4253 = i == 8'h0 ? _GEN_4252 : _GEN_2863; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4254 = io_inputBit | _GEN_4253; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4255 = i == 8'h2 ? _GEN_4254 : _GEN_4253; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4256 = io_inputBit | _GEN_4255; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4257 = i == 8'h5 ? _GEN_4256 : _GEN_4255; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4258 = io_inputBit | _GEN_4257; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4259 = i == 8'hb ? _GEN_4258 : _GEN_4257; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4260 = ~io_inputBit ? 1'h0 : _GEN_4259; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4261 = i == 8'h17 ? _GEN_4260 : _GEN_4259; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4262 = ~io_inputBit ? 1'h0 : _GEN_4261; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4263 = i == 8'h30 ? _GEN_4262 : _GEN_4261; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4264 = io_inputBit | _GEN_4263; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4265 = i == 8'h62 ? _GEN_4264 : _GEN_4263; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4266 = ~io_inputBit ? 1'h0 : _GEN_4265; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4267 = i == 8'hc5 ? _GEN_4266 : _GEN_4265; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4268 = io_inputBit | _GEN_4267; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4269 = i == 8'hc5 ? _GEN_4268 : _GEN_4267; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4270 = ~io_inputBit ? 1'h0 : _GEN_2943; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4271 = i == 8'h0 ? _GEN_4270 : _GEN_2943; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4272 = io_inputBit | _GEN_4271; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4273 = i == 8'h2 ? _GEN_4272 : _GEN_4271; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4274 = io_inputBit | _GEN_4273; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4275 = i == 8'h5 ? _GEN_4274 : _GEN_4273; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4276 = io_inputBit | _GEN_4275; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4277 = i == 8'h18 ? _GEN_4276 : _GEN_4275; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4278 = ~io_inputBit ? 1'h0 : _GEN_4277; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4279 = i == 8'h2f ? _GEN_4278 : _GEN_4277; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4280 = ~io_inputBit | _GEN_4279; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4281 = i == 8'h30 ? _GEN_4280 : _GEN_4279; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4282 = ~io_inputBit ? 1'h0 : _GEN_4281; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4283 = i == 8'h31 ? _GEN_4282 : _GEN_4281; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4284 = io_inputBit | _GEN_4283; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4285 = i == 8'h60 ? _GEN_4284 : _GEN_4283; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4286 = io_inputBit ? 1'h0 : _GEN_4285; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4287 = i == 8'h62 ? _GEN_4286 : _GEN_4285; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4288 = io_inputBit | _GEN_4287; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4289 = i == 8'h64 ? _GEN_4288 : _GEN_4287; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4290 = ~io_inputBit ? 1'h0 : _GEN_4289; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4291 = i == 8'hc1 ? _GEN_4290 : _GEN_4289; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4292 = io_inputBit | _GEN_4291; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4293 = i == 8'hc1 ? _GEN_4292 : _GEN_4291; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4294 = ~io_inputBit | _GEN_4293; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4295 = i == 8'hc5 ? _GEN_4294 : _GEN_4293; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4296 = io_inputBit ? 1'h0 : _GEN_4295; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4297 = i == 8'hc5 ? _GEN_4296 : _GEN_4295; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4298 = ~io_inputBit ? 1'h0 : _GEN_4297; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4299 = i == 8'hc9 ? _GEN_4298 : _GEN_4297; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4300 = io_inputBit | _GEN_4299; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4301 = i == 8'hc9 ? _GEN_4300 : _GEN_4299; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4302 = ~io_inputBit ? 1'h0 : _GEN_3065; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4303 = i == 8'h0 ? _GEN_4302 : _GEN_3065; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4304 = io_inputBit ? 1'h0 : _GEN_4303; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4305 = i == 8'h2 ? _GEN_4304 : _GEN_4303; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4306 = io_inputBit ? 1'h0 : _GEN_4305; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4307 = i == 8'h5 ? _GEN_4306 : _GEN_4305; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4308 = io_inputBit ? 1'h0 : _GEN_4307; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4309 = i == 8'h18 ? _GEN_4308 : _GEN_4307; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4310 = io_inputBit | _GEN_4309; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4311 = i == 8'h5f ? _GEN_4310 : _GEN_4309; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4312 = io_inputBit ? 1'h0 : _GEN_4311; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4313 = i == 8'h60 ? _GEN_4312 : _GEN_4311; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4314 = io_inputBit | _GEN_4313; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4315 = i == 8'h61 ? _GEN_4314 : _GEN_4313; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4316 = io_inputBit ? 1'h0 : _GEN_4315; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4317 = i == 8'h62 ? _GEN_4316 : _GEN_4315; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4318 = io_inputBit | _GEN_4317; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4319 = i == 8'h63 ? _GEN_4318 : _GEN_4317; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4320 = io_inputBit ? 1'h0 : _GEN_4319; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4321 = i == 8'h64 ? _GEN_4320 : _GEN_4319; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4322 = ~io_inputBit ? 1'h0 : _GEN_4321; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4323 = i == 8'hbf ? _GEN_4322 : _GEN_4321; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4324 = io_inputBit | _GEN_4323; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4325 = i == 8'hbf ? _GEN_4324 : _GEN_4323; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4326 = ~io_inputBit | _GEN_4325; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4327 = i == 8'hc1 ? _GEN_4326 : _GEN_4325; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4328 = io_inputBit ? 1'h0 : _GEN_4327; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4329 = i == 8'hc1 ? _GEN_4328 : _GEN_4327; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4330 = ~io_inputBit ? 1'h0 : _GEN_4329; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4331 = i == 8'hc3 ? _GEN_4330 : _GEN_4329; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4332 = io_inputBit | _GEN_4331; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4333 = i == 8'hc3 ? _GEN_4332 : _GEN_4331; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4334 = ~io_inputBit | _GEN_4333; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4335 = i == 8'hc5 ? _GEN_4334 : _GEN_4333; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4336 = io_inputBit ? 1'h0 : _GEN_4335; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4337 = i == 8'hc5 ? _GEN_4336 : _GEN_4335; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4338 = ~io_inputBit ? 1'h0 : _GEN_4337; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4339 = i == 8'hc7 ? _GEN_4338 : _GEN_4337; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4340 = io_inputBit | _GEN_4339; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4341 = i == 8'hc7 ? _GEN_4340 : _GEN_4339; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4342 = ~io_inputBit | _GEN_4341; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4343 = i == 8'hc9 ? _GEN_4342 : _GEN_4341; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4344 = io_inputBit ? 1'h0 : _GEN_4343; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4345 = i == 8'hc9 ? _GEN_4344 : _GEN_4343; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4346 = ~io_inputBit ? 1'h0 : _GEN_3247; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4347 = i == 8'h1 ? _GEN_4346 : _GEN_3247; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4348 = io_inputBit ? 1'h0 : _GEN_4347; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4349 = i == 8'h2 ? _GEN_4348 : _GEN_4347; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4350 = ~io_inputBit ? 1'h0 : _GEN_4349; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4351 = i == 8'h4 ? _GEN_4350 : _GEN_4349; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4352 = io_inputBit ? 1'h0 : _GEN_4351; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4353 = i == 8'h5 ? _GEN_4352 : _GEN_4351; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4354 = ~io_inputBit ? 1'h0 : _GEN_4353; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4355 = i == 8'ha ? _GEN_4354 : _GEN_4353; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4356 = ~io_inputBit ? 1'h0 : _GEN_4355; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4357 = i == 8'h16 ? _GEN_4356 : _GEN_4355; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4358 = io_inputBit ? 1'h0 : _GEN_4357; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4359 = i == 8'h18 ? _GEN_4358 : _GEN_4357; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4360 = ~io_inputBit ? 1'h0 : _GEN_4359; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4361 = i == 8'h2e ? _GEN_4360 : _GEN_4359; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4362 = ~io_inputBit ? 1'h0 : _GEN_4361; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4363 = i == 8'h5e ? _GEN_4362 : _GEN_4361; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4364 = io_inputBit ? 1'h0 : _GEN_4363; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4365 = i == 8'h64 ? _GEN_4364 : _GEN_4363; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4366 = ~io_inputBit ? 1'h0 : _GEN_4365; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4367 = i == 8'hbe ? _GEN_4366 : _GEN_4365; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4368 = io_inputBit | _GEN_4367; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4369 = i == 8'hbe ? _GEN_4368 : _GEN_4367; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4370 = ~io_inputBit | _GEN_4369; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4371 = i == 8'hbf ? _GEN_4370 : _GEN_4369; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4372 = io_inputBit ? 1'h0 : _GEN_4371; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4373 = i == 8'hbf ? _GEN_4372 : _GEN_4371; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4374 = ~io_inputBit ? 1'h0 : _GEN_4373; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4375 = i == 8'hc0 ? _GEN_4374 : _GEN_4373; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4376 = io_inputBit | _GEN_4375; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4377 = i == 8'hc0 ? _GEN_4376 : _GEN_4375; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4378 = ~io_inputBit | _GEN_4377; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4379 = i == 8'hc1 ? _GEN_4378 : _GEN_4377; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4380 = io_inputBit ? 1'h0 : _GEN_4379; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4381 = i == 8'hc1 ? _GEN_4380 : _GEN_4379; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4382 = ~io_inputBit ? 1'h0 : _GEN_4381; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4383 = i == 8'hc2 ? _GEN_4382 : _GEN_4381; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4384 = io_inputBit | _GEN_4383; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4385 = i == 8'hc2 ? _GEN_4384 : _GEN_4383; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4386 = ~io_inputBit | _GEN_4385; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4387 = i == 8'hc3 ? _GEN_4386 : _GEN_4385; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4388 = io_inputBit ? 1'h0 : _GEN_4387; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4389 = i == 8'hc3 ? _GEN_4388 : _GEN_4387; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4390 = ~io_inputBit ? 1'h0 : _GEN_4389; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4391 = i == 8'hc4 ? _GEN_4390 : _GEN_4389; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4392 = io_inputBit | _GEN_4391; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4393 = i == 8'hc4 ? _GEN_4392 : _GEN_4391; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4394 = ~io_inputBit | _GEN_4393; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4395 = i == 8'hc5 ? _GEN_4394 : _GEN_4393; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4396 = io_inputBit ? 1'h0 : _GEN_4395; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4397 = i == 8'hc5 ? _GEN_4396 : _GEN_4395; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4398 = ~io_inputBit ? 1'h0 : _GEN_4397; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4399 = i == 8'hc6 ? _GEN_4398 : _GEN_4397; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4400 = io_inputBit | _GEN_4399; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4401 = i == 8'hc6 ? _GEN_4400 : _GEN_4399; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4402 = ~io_inputBit | _GEN_4401; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4403 = i == 8'hc7 ? _GEN_4402 : _GEN_4401; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4404 = io_inputBit ? 1'h0 : _GEN_4403; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4405 = i == 8'hc7 ? _GEN_4404 : _GEN_4403; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4406 = ~io_inputBit ? 1'h0 : _GEN_4405; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4407 = i == 8'hc8 ? _GEN_4406 : _GEN_4405; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4408 = io_inputBit | _GEN_4407; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4409 = i == 8'hc8 ? _GEN_4408 : _GEN_4407; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4410 = ~io_inputBit | _GEN_4409; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4411 = i == 8'hc9 ? _GEN_4410 : _GEN_4409; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4412 = io_inputBit ? 1'h0 : _GEN_4411; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4413 = i == 8'hc9 ? _GEN_4412 : _GEN_4411; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4414 = ~io_inputBit ? 1'h0 : _GEN_3511; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4415 = i == 8'h1 ? _GEN_4414 : _GEN_3511; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4416 = io_inputBit | _GEN_4415; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4417 = i == 8'h2 ? _GEN_4416 : _GEN_4415; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4418 = ~io_inputBit ? 1'h0 : _GEN_4417; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4419 = i == 8'h4 ? _GEN_4418 : _GEN_4417; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4420 = io_inputBit | _GEN_4419; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4421 = i == 8'h5 ? _GEN_4420 : _GEN_4419; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4422 = ~io_inputBit ? 1'h0 : _GEN_4421; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4423 = i == 8'ha ? _GEN_4422 : _GEN_4421; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4424 = ~io_inputBit ? 1'h0 : _GEN_4423; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4425 = i == 8'h16 ? _GEN_4424 : _GEN_4423; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4426 = io_inputBit | _GEN_4425; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4427 = i == 8'h18 ? _GEN_4426 : _GEN_4425; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4428 = ~io_inputBit ? 1'h0 : _GEN_4427; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4429 = i == 8'h2e ? _GEN_4428 : _GEN_4427; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4430 = ~io_inputBit ? 1'h0 : _GEN_4429; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4431 = i == 8'h5e ? _GEN_4430 : _GEN_4429; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4432 = io_inputBit | _GEN_4431; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4433 = i == 8'h64 ? _GEN_4432 : _GEN_4431; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4434 = ~io_inputBit | _GEN_4433; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4435 = i == 8'hbe ? _GEN_4434 : _GEN_4433; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4436 = io_inputBit ? 1'h0 : _GEN_4435; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4437 = i == 8'hbe ? _GEN_4436 : _GEN_4435; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4438 = ~io_inputBit | _GEN_4437; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4439 = i == 8'hbf ? _GEN_4438 : _GEN_4437; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4440 = io_inputBit ? 1'h0 : _GEN_4439; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4441 = i == 8'hbf ? _GEN_4440 : _GEN_4439; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4442 = ~io_inputBit | _GEN_4441; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4443 = i == 8'hc0 ? _GEN_4442 : _GEN_4441; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4444 = io_inputBit ? 1'h0 : _GEN_4443; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4445 = i == 8'hc0 ? _GEN_4444 : _GEN_4443; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4446 = ~io_inputBit | _GEN_4445; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4447 = i == 8'hc1 ? _GEN_4446 : _GEN_4445; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4448 = io_inputBit ? 1'h0 : _GEN_4447; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4449 = i == 8'hc1 ? _GEN_4448 : _GEN_4447; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4450 = ~io_inputBit | _GEN_4449; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4451 = i == 8'hc2 ? _GEN_4450 : _GEN_4449; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4452 = io_inputBit ? 1'h0 : _GEN_4451; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4453 = i == 8'hc2 ? _GEN_4452 : _GEN_4451; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4454 = ~io_inputBit | _GEN_4453; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4455 = i == 8'hc3 ? _GEN_4454 : _GEN_4453; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4456 = io_inputBit ? 1'h0 : _GEN_4455; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4457 = i == 8'hc3 ? _GEN_4456 : _GEN_4455; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4458 = ~io_inputBit | _GEN_4457; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4459 = i == 8'hc4 ? _GEN_4458 : _GEN_4457; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4460 = io_inputBit ? 1'h0 : _GEN_4459; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4461 = i == 8'hc4 ? _GEN_4460 : _GEN_4459; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4462 = ~io_inputBit | _GEN_4461; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4463 = i == 8'hc5 ? _GEN_4462 : _GEN_4461; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4464 = io_inputBit ? 1'h0 : _GEN_4463; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4465 = i == 8'hc5 ? _GEN_4464 : _GEN_4463; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4466 = ~io_inputBit | _GEN_4465; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4467 = i == 8'hc6 ? _GEN_4466 : _GEN_4465; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4468 = io_inputBit ? 1'h0 : _GEN_4467; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4469 = i == 8'hc6 ? _GEN_4468 : _GEN_4467; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4470 = ~io_inputBit | _GEN_4469; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4471 = i == 8'hc7 ? _GEN_4470 : _GEN_4469; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4472 = io_inputBit ? 1'h0 : _GEN_4471; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4473 = i == 8'hc7 ? _GEN_4472 : _GEN_4471; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4474 = ~io_inputBit | _GEN_4473; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4475 = i == 8'hc8 ? _GEN_4474 : _GEN_4473; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4476 = io_inputBit ? 1'h0 : _GEN_4475; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4477 = i == 8'hc8 ? _GEN_4476 : _GEN_4475; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4478 = ~io_inputBit | _GEN_4477; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4479 = i == 8'hc9 ? _GEN_4478 : _GEN_4477; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4480 = io_inputBit ? 1'h0 : _GEN_4479; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4481 = i == 8'hc9 ? _GEN_4480 : _GEN_4479; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4482 = ~io_inputBit ? 1'h0 : _GEN_3827; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4483 = i == 8'h1 ? _GEN_4482 : _GEN_3827; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4484 = io_inputBit ? 1'h0 : _GEN_4483; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4485 = i == 8'h2 ? _GEN_4484 : _GEN_4483; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4486 = ~io_inputBit ? 1'h0 : _GEN_4485; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4487 = i == 8'h4 ? _GEN_4486 : _GEN_4485; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4488 = io_inputBit ? 1'h0 : _GEN_4487; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4489 = i == 8'h5 ? _GEN_4488 : _GEN_4487; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4490 = ~io_inputBit ? 1'h0 : _GEN_4489; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4491 = i == 8'ha ? _GEN_4490 : _GEN_4489; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4492 = ~io_inputBit ? 1'h0 : _GEN_4491; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4493 = i == 8'h16 ? _GEN_4492 : _GEN_4491; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4494 = io_inputBit ? 1'h0 : _GEN_4493; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4495 = i == 8'h18 ? _GEN_4494 : _GEN_4493; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4496 = ~io_inputBit ? 1'h0 : _GEN_4495; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4497 = i == 8'h2e ? _GEN_4496 : _GEN_4495; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4498 = io_inputBit ? 1'h0 : _GEN_4497; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4499 = i == 8'h64 ? _GEN_4498 : _GEN_4497; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4500 = ~io_inputBit ? 1'h0 : _GEN_4499; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4501 = i == 8'hbd ? _GEN_4500 : _GEN_4499; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4502 = ~io_inputBit ? 1'h0 : _GEN_4501; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4503 = _GEN_6084 == 9'h17c ? _GEN_4502 : _GEN_4501; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4504 = io_inputBit | _GEN_4503; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4505 = _GEN_6084 == 9'h17c ? _GEN_4504 : _GEN_4503; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4506 = ~io_inputBit ? 1'h0 : _GEN_4505; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4507 = _GEN_6084 == 9'h17d ? _GEN_4506 : _GEN_4505; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4508 = io_inputBit | _GEN_4507; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4509 = _GEN_6084 == 9'h17d ? _GEN_4508 : _GEN_4507; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4510 = ~io_inputBit ? 1'h0 : _GEN_4509; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4511 = _GEN_6084 == 9'h17e ? _GEN_4510 : _GEN_4509; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4512 = io_inputBit | _GEN_4511; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4513 = _GEN_6084 == 9'h17e ? _GEN_4512 : _GEN_4511; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4514 = ~io_inputBit ? 1'h0 : _GEN_4513; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4515 = _GEN_6084 == 9'h17f ? _GEN_4514 : _GEN_4513; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4516 = io_inputBit | _GEN_4515; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4517 = _GEN_6084 == 9'h17f ? _GEN_4516 : _GEN_4515; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4518 = ~io_inputBit ? 1'h0 : _GEN_4517; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4519 = _GEN_6084 == 9'h180 ? _GEN_4518 : _GEN_4517; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4520 = io_inputBit | _GEN_4519; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4521 = _GEN_6084 == 9'h180 ? _GEN_4520 : _GEN_4519; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4522 = ~io_inputBit ? 1'h0 : _GEN_4521; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4523 = _GEN_6084 == 9'h181 ? _GEN_4522 : _GEN_4521; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4524 = io_inputBit | _GEN_4523; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4525 = _GEN_6084 == 9'h181 ? _GEN_4524 : _GEN_4523; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4526 = ~io_inputBit ? 1'h0 : _GEN_4525; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4527 = _GEN_6084 == 9'h182 ? _GEN_4526 : _GEN_4525; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4528 = io_inputBit | _GEN_4527; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4529 = _GEN_6084 == 9'h182 ? _GEN_4528 : _GEN_4527; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4530 = ~io_inputBit ? 1'h0 : _GEN_4529; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4531 = _GEN_6084 == 9'h183 ? _GEN_4530 : _GEN_4529; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4532 = io_inputBit | _GEN_4531; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4533 = _GEN_6084 == 9'h183 ? _GEN_4532 : _GEN_4531; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4534 = ~io_inputBit ? 1'h0 : _GEN_4533; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4535 = _GEN_6084 == 9'h184 ? _GEN_4534 : _GEN_4533; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4536 = io_inputBit | _GEN_4535; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4537 = _GEN_6084 == 9'h184 ? _GEN_4536 : _GEN_4535; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4538 = ~io_inputBit ? 1'h0 : _GEN_4537; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4539 = _GEN_6084 == 9'h185 ? _GEN_4538 : _GEN_4537; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4540 = io_inputBit | _GEN_4539; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4541 = _GEN_6084 == 9'h185 ? _GEN_4540 : _GEN_4539; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4542 = ~io_inputBit ? 1'h0 : _GEN_4541; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4543 = _GEN_6084 == 9'h186 ? _GEN_4542 : _GEN_4541; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4544 = io_inputBit | _GEN_4543; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4545 = _GEN_6084 == 9'h186 ? _GEN_4544 : _GEN_4543; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4546 = ~io_inputBit ? 1'h0 : _GEN_4545; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4547 = _GEN_6084 == 9'h187 ? _GEN_4546 : _GEN_4545; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4548 = io_inputBit | _GEN_4547; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4549 = _GEN_6084 == 9'h187 ? _GEN_4548 : _GEN_4547; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4550 = ~io_inputBit ? 1'h0 : _GEN_4549; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4551 = _GEN_6084 == 9'h188 ? _GEN_4550 : _GEN_4549; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4552 = io_inputBit | _GEN_4551; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4553 = _GEN_6084 == 9'h188 ? _GEN_4552 : _GEN_4551; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4554 = ~io_inputBit ? 1'h0 : _GEN_4553; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4555 = _GEN_6084 == 9'h189 ? _GEN_4554 : _GEN_4553; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4556 = io_inputBit | _GEN_4555; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4557 = _GEN_6084 == 9'h189 ? _GEN_4556 : _GEN_4555; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4558 = ~io_inputBit ? 1'h0 : _GEN_4557; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4559 = _GEN_6084 == 9'h18a ? _GEN_4558 : _GEN_4557; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4560 = io_inputBit | _GEN_4559; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4561 = _GEN_6084 == 9'h18a ? _GEN_4560 : _GEN_4559; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4562 = ~io_inputBit ? 1'h0 : _GEN_4561; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4563 = _GEN_6084 == 9'h18b ? _GEN_4562 : _GEN_4561; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4564 = io_inputBit | _GEN_4563; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4565 = _GEN_6084 == 9'h18b ? _GEN_4564 : _GEN_4563; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4566 = ~io_inputBit ? 1'h0 : _GEN_4565; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4567 = _GEN_6084 == 9'h18c ? _GEN_4566 : _GEN_4565; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4568 = io_inputBit | _GEN_4567; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4569 = _GEN_6084 == 9'h18c ? _GEN_4568 : _GEN_4567; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4570 = ~io_inputBit ? 1'h0 : _GEN_4569; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4571 = _GEN_6084 == 9'h18d ? _GEN_4570 : _GEN_4569; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4572 = io_inputBit | _GEN_4571; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4573 = _GEN_6084 == 9'h18d ? _GEN_4572 : _GEN_4571; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4574 = ~io_inputBit ? 1'h0 : _GEN_4573; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4575 = _GEN_6084 == 9'h18e ? _GEN_4574 : _GEN_4573; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4576 = io_inputBit | _GEN_4575; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4577 = _GEN_6084 == 9'h18e ? _GEN_4576 : _GEN_4575; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4578 = ~io_inputBit ? 1'h0 : _GEN_4577; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4579 = _GEN_6084 == 9'h18f ? _GEN_4578 : _GEN_4577; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4580 = io_inputBit | _GEN_4579; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4581 = _GEN_6084 == 9'h18f ? _GEN_4580 : _GEN_4579; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4582 = ~io_inputBit ? 1'h0 : _GEN_4581; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4583 = _GEN_6084 == 9'h190 ? _GEN_4582 : _GEN_4581; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4584 = io_inputBit | _GEN_4583; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4585 = _GEN_6084 == 9'h190 ? _GEN_4584 : _GEN_4583; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4586 = ~io_inputBit ? 1'h0 : _GEN_4585; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4587 = _GEN_6084 == 9'h191 ? _GEN_4586 : _GEN_4585; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4588 = io_inputBit | _GEN_4587; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4589 = _GEN_6084 == 9'h191 ? _GEN_4588 : _GEN_4587; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4590 = ~io_inputBit ? 1'h0 : _GEN_4589; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4591 = _GEN_6084 == 9'h192 ? _GEN_4590 : _GEN_4589; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4592 = io_inputBit | _GEN_4591; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4593 = _GEN_6084 == 9'h192 ? _GEN_4592 : _GEN_4591; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4594 = ~io_inputBit ? 1'h0 : _GEN_4593; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4595 = _GEN_6084 == 9'h193 ? _GEN_4594 : _GEN_4593; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4596 = io_inputBit | _GEN_4595; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4597 = _GEN_6084 == 9'h193 ? _GEN_4596 : _GEN_4595; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4598 = ~io_inputBit ? 1'h0 : _GEN_4597; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4599 = _GEN_6084 == 9'h194 ? _GEN_4598 : _GEN_4597; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4600 = io_inputBit | _GEN_4599; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4601 = _GEN_6084 == 9'h194 ? _GEN_4600 : _GEN_4599; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4602 = ~io_inputBit ? 1'h0 : _GEN_4251; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4603 = i == 8'h1 ? _GEN_4602 : _GEN_4251; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4604 = io_inputBit ? 1'h0 : _GEN_4603; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4605 = i == 8'h2 ? _GEN_4604 : _GEN_4603; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4606 = ~io_inputBit ? 1'h0 : _GEN_4605; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4607 = i == 8'h4 ? _GEN_4606 : _GEN_4605; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4608 = io_inputBit ? 1'h0 : _GEN_4607; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4609 = i == 8'h5 ? _GEN_4608 : _GEN_4607; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4610 = ~io_inputBit ? 1'h0 : _GEN_4609; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4611 = i == 8'ha ? _GEN_4610 : _GEN_4609; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4612 = ~io_inputBit ? 1'h0 : _GEN_4611; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4613 = i == 8'h16 ? _GEN_4612 : _GEN_4611; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4614 = io_inputBit ? 1'h0 : _GEN_4613; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4615 = i == 8'h18 ? _GEN_4614 : _GEN_4613; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4616 = ~io_inputBit ? 1'h0 : _GEN_4615; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4617 = i == 8'h2e ? _GEN_4616 : _GEN_4615; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4618 = io_inputBit ? 1'h0 : _GEN_4617; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4619 = i == 8'h64 ? _GEN_4618 : _GEN_4617; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4620 = ~io_inputBit ? 1'h0 : _GEN_4619; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4621 = i == 8'hbd ? _GEN_4620 : _GEN_4619; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4622 = ~io_inputBit ? 1'h0 : _GEN_4621; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4623 = _GEN_6085 == 10'h2f9 ? _GEN_4622 : _GEN_4621; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4624 = io_inputBit | _GEN_4623; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4625 = _GEN_6085 == 10'h2f9 ? _GEN_4624 : _GEN_4623; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4626 = ~io_inputBit ? 1'h0 : _GEN_4625; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4627 = _GEN_6085 == 10'h2fa ? _GEN_4626 : _GEN_4625; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4628 = io_inputBit | _GEN_4627; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4629 = _GEN_6085 == 10'h2fa ? _GEN_4628 : _GEN_4627; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4630 = ~io_inputBit ? 1'h0 : _GEN_4629; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4631 = _GEN_6085 == 10'h2fb ? _GEN_4630 : _GEN_4629; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4632 = io_inputBit | _GEN_4631; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4633 = _GEN_6085 == 10'h2fb ? _GEN_4632 : _GEN_4631; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4634 = ~io_inputBit ? 1'h0 : _GEN_4633; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4635 = _GEN_6085 == 10'h2fc ? _GEN_4634 : _GEN_4633; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4636 = io_inputBit | _GEN_4635; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4637 = _GEN_6085 == 10'h2fc ? _GEN_4636 : _GEN_4635; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4638 = ~io_inputBit ? 1'h0 : _GEN_4637; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4639 = _GEN_6085 == 10'h2fd ? _GEN_4638 : _GEN_4637; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4640 = io_inputBit | _GEN_4639; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4641 = _GEN_6085 == 10'h2fd ? _GEN_4640 : _GEN_4639; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4642 = ~io_inputBit ? 1'h0 : _GEN_4641; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4643 = _GEN_6085 == 10'h2fe ? _GEN_4642 : _GEN_4641; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4644 = io_inputBit | _GEN_4643; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4645 = _GEN_6085 == 10'h2fe ? _GEN_4644 : _GEN_4643; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4646 = ~io_inputBit ? 1'h0 : _GEN_4645; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4647 = _GEN_6085 == 10'h2ff ? _GEN_4646 : _GEN_4645; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4648 = io_inputBit | _GEN_4647; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4649 = _GEN_6085 == 10'h2ff ? _GEN_4648 : _GEN_4647; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4650 = ~io_inputBit ? 1'h0 : _GEN_4649; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4651 = _GEN_6085 == 10'h300 ? _GEN_4650 : _GEN_4649; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4652 = io_inputBit | _GEN_4651; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4653 = _GEN_6085 == 10'h300 ? _GEN_4652 : _GEN_4651; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4654 = ~io_inputBit ? 1'h0 : _GEN_4653; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4655 = _GEN_6085 == 10'h301 ? _GEN_4654 : _GEN_4653; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4656 = io_inputBit | _GEN_4655; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4657 = _GEN_6085 == 10'h301 ? _GEN_4656 : _GEN_4655; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4658 = ~io_inputBit ? 1'h0 : _GEN_4657; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4659 = _GEN_6085 == 10'h302 ? _GEN_4658 : _GEN_4657; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4660 = io_inputBit | _GEN_4659; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4661 = _GEN_6085 == 10'h302 ? _GEN_4660 : _GEN_4659; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4662 = ~io_inputBit ? 1'h0 : _GEN_4661; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4663 = _GEN_6085 == 10'h303 ? _GEN_4662 : _GEN_4661; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4664 = io_inputBit | _GEN_4663; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4665 = _GEN_6085 == 10'h303 ? _GEN_4664 : _GEN_4663; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4666 = ~io_inputBit ? 1'h0 : _GEN_4665; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4667 = _GEN_6085 == 10'h304 ? _GEN_4666 : _GEN_4665; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4668 = io_inputBit | _GEN_4667; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4669 = _GEN_6085 == 10'h304 ? _GEN_4668 : _GEN_4667; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4670 = ~io_inputBit ? 1'h0 : _GEN_4669; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4671 = _GEN_6085 == 10'h305 ? _GEN_4670 : _GEN_4669; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4672 = io_inputBit | _GEN_4671; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4673 = _GEN_6085 == 10'h305 ? _GEN_4672 : _GEN_4671; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4674 = ~io_inputBit ? 1'h0 : _GEN_4673; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4675 = _GEN_6085 == 10'h306 ? _GEN_4674 : _GEN_4673; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4676 = io_inputBit | _GEN_4675; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4677 = _GEN_6085 == 10'h306 ? _GEN_4676 : _GEN_4675; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4678 = ~io_inputBit ? 1'h0 : _GEN_4677; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4679 = _GEN_6085 == 10'h307 ? _GEN_4678 : _GEN_4677; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4680 = io_inputBit | _GEN_4679; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4681 = _GEN_6085 == 10'h307 ? _GEN_4680 : _GEN_4679; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4682 = ~io_inputBit ? 1'h0 : _GEN_4681; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4683 = _GEN_6085 == 10'h308 ? _GEN_4682 : _GEN_4681; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4684 = io_inputBit | _GEN_4683; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4685 = _GEN_6085 == 10'h308 ? _GEN_4684 : _GEN_4683; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4686 = ~io_inputBit ? 1'h0 : _GEN_4685; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4687 = _GEN_6085 == 10'h309 ? _GEN_4686 : _GEN_4685; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4688 = io_inputBit | _GEN_4687; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4689 = _GEN_6085 == 10'h309 ? _GEN_4688 : _GEN_4687; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4690 = ~io_inputBit ? 1'h0 : _GEN_4689; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4691 = _GEN_6085 == 10'h30a ? _GEN_4690 : _GEN_4689; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4692 = io_inputBit | _GEN_4691; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4693 = _GEN_6085 == 10'h30a ? _GEN_4692 : _GEN_4691; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4694 = ~io_inputBit ? 1'h0 : _GEN_4693; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4695 = _GEN_6085 == 10'h30b ? _GEN_4694 : _GEN_4693; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4696 = io_inputBit | _GEN_4695; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4697 = _GEN_6085 == 10'h30b ? _GEN_4696 : _GEN_4695; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4698 = ~io_inputBit ? 1'h0 : _GEN_4697; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4699 = _GEN_6085 == 10'h30c ? _GEN_4698 : _GEN_4697; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4700 = io_inputBit | _GEN_4699; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4701 = _GEN_6085 == 10'h30c ? _GEN_4700 : _GEN_4699; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4702 = ~io_inputBit ? 1'h0 : _GEN_4701; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4703 = _GEN_6085 == 10'h30d ? _GEN_4702 : _GEN_4701; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4704 = io_inputBit | _GEN_4703; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4705 = _GEN_6085 == 10'h30d ? _GEN_4704 : _GEN_4703; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4706 = ~io_inputBit ? 1'h0 : _GEN_4705; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4707 = _GEN_6085 == 10'h30e ? _GEN_4706 : _GEN_4705; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4708 = io_inputBit | _GEN_4707; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4709 = _GEN_6085 == 10'h30e ? _GEN_4708 : _GEN_4707; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4710 = ~io_inputBit ? 1'h0 : _GEN_4709; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4711 = _GEN_6085 == 10'h30f ? _GEN_4710 : _GEN_4709; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4712 = io_inputBit | _GEN_4711; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4713 = _GEN_6085 == 10'h30f ? _GEN_4712 : _GEN_4711; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4714 = ~io_inputBit ? 1'h0 : _GEN_4713; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4715 = _GEN_6085 == 10'h310 ? _GEN_4714 : _GEN_4713; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4716 = io_inputBit | _GEN_4715; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4717 = _GEN_6085 == 10'h310 ? _GEN_4716 : _GEN_4715; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4718 = ~io_inputBit ? 1'h0 : _GEN_4717; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4719 = _GEN_6085 == 10'h311 ? _GEN_4718 : _GEN_4717; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4720 = io_inputBit | _GEN_4719; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4721 = _GEN_6085 == 10'h311 ? _GEN_4720 : _GEN_4719; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4722 = ~io_inputBit ? 1'h0 : _GEN_4721; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4723 = _GEN_6085 == 10'h312 ? _GEN_4722 : _GEN_4721; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4724 = io_inputBit | _GEN_4723; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4725 = _GEN_6085 == 10'h312 ? _GEN_4724 : _GEN_4723; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4726 = ~io_inputBit ? 1'h0 : _GEN_4725; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4727 = _GEN_6085 == 10'h313 ? _GEN_4726 : _GEN_4725; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4728 = io_inputBit | _GEN_4727; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4729 = _GEN_6085 == 10'h313 ? _GEN_4728 : _GEN_4727; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4730 = ~io_inputBit ? 1'h0 : _GEN_4729; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4731 = _GEN_6085 == 10'h314 ? _GEN_4730 : _GEN_4729; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4732 = io_inputBit | _GEN_4731; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4733 = _GEN_6085 == 10'h314 ? _GEN_4732 : _GEN_4731; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4734 = ~io_inputBit ? 1'h0 : _GEN_4733; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4735 = _GEN_6085 == 10'h315 ? _GEN_4734 : _GEN_4733; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4736 = io_inputBit | _GEN_4735; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4737 = _GEN_6085 == 10'h315 ? _GEN_4736 : _GEN_4735; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4738 = ~io_inputBit ? 1'h0 : _GEN_4737; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4739 = _GEN_6085 == 10'h316 ? _GEN_4738 : _GEN_4737; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4740 = io_inputBit | _GEN_4739; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4741 = _GEN_6085 == 10'h316 ? _GEN_4740 : _GEN_4739; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4742 = ~io_inputBit ? 1'h0 : _GEN_4741; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4743 = _GEN_6085 == 10'h317 ? _GEN_4742 : _GEN_4741; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4744 = io_inputBit | _GEN_4743; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4745 = _GEN_6085 == 10'h317 ? _GEN_4744 : _GEN_4743; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4746 = ~io_inputBit ? 1'h0 : _GEN_4745; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4747 = _GEN_6085 == 10'h318 ? _GEN_4746 : _GEN_4745; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4748 = io_inputBit | _GEN_4747; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4749 = _GEN_6085 == 10'h318 ? _GEN_4748 : _GEN_4747; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4750 = ~io_inputBit ? 1'h0 : _GEN_4749; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4751 = _GEN_6085 == 10'h319 ? _GEN_4750 : _GEN_4749; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4752 = io_inputBit | _GEN_4751; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4753 = _GEN_6085 == 10'h319 ? _GEN_4752 : _GEN_4751; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4754 = ~io_inputBit ? 1'h0 : _GEN_4753; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4755 = _GEN_6085 == 10'h31a ? _GEN_4754 : _GEN_4753; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4756 = io_inputBit | _GEN_4755; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4757 = _GEN_6085 == 10'h31a ? _GEN_4756 : _GEN_4755; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4758 = ~io_inputBit ? 1'h0 : _GEN_4757; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4759 = _GEN_6085 == 10'h31b ? _GEN_4758 : _GEN_4757; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4760 = io_inputBit | _GEN_4759; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4761 = _GEN_6085 == 10'h31b ? _GEN_4760 : _GEN_4759; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4762 = ~io_inputBit ? 1'h0 : _GEN_4761; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4763 = _GEN_6085 == 10'h31c ? _GEN_4762 : _GEN_4761; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4764 = io_inputBit | _GEN_4763; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4765 = _GEN_6085 == 10'h31c ? _GEN_4764 : _GEN_4763; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4766 = ~io_inputBit ? 1'h0 : _GEN_4765; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4767 = _GEN_6085 == 10'h31d ? _GEN_4766 : _GEN_4765; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4768 = io_inputBit | _GEN_4767; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4769 = _GEN_6085 == 10'h31d ? _GEN_4768 : _GEN_4767; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4770 = ~io_inputBit ? 1'h0 : _GEN_4769; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4771 = _GEN_6085 == 10'h31e ? _GEN_4770 : _GEN_4769; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4772 = io_inputBit | _GEN_4771; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4773 = _GEN_6085 == 10'h31e ? _GEN_4772 : _GEN_4771; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4774 = ~io_inputBit ? 1'h0 : _GEN_4773; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4775 = _GEN_6085 == 10'h31f ? _GEN_4774 : _GEN_4773; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4776 = io_inputBit | _GEN_4775; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4777 = _GEN_6085 == 10'h31f ? _GEN_4776 : _GEN_4775; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4778 = ~io_inputBit ? 1'h0 : _GEN_4777; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4779 = _GEN_6085 == 10'h320 ? _GEN_4778 : _GEN_4777; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4780 = io_inputBit | _GEN_4779; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4781 = _GEN_6085 == 10'h320 ? _GEN_4780 : _GEN_4779; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4782 = ~io_inputBit ? 1'h0 : _GEN_4781; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4783 = _GEN_6085 == 10'h321 ? _GEN_4782 : _GEN_4781; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4784 = io_inputBit | _GEN_4783; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4785 = _GEN_6085 == 10'h321 ? _GEN_4784 : _GEN_4783; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4786 = ~io_inputBit ? 1'h0 : _GEN_4785; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4787 = _GEN_6085 == 10'h322 ? _GEN_4786 : _GEN_4785; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4788 = io_inputBit | _GEN_4787; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4789 = _GEN_6085 == 10'h322 ? _GEN_4788 : _GEN_4787; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4790 = ~io_inputBit ? 1'h0 : _GEN_4789; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4791 = _GEN_6085 == 10'h323 ? _GEN_4790 : _GEN_4789; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4792 = io_inputBit | _GEN_4791; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4793 = _GEN_6085 == 10'h323 ? _GEN_4792 : _GEN_4791; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4794 = ~io_inputBit ? 1'h0 : _GEN_4793; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4795 = _GEN_6085 == 10'h324 ? _GEN_4794 : _GEN_4793; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4796 = io_inputBit | _GEN_4795; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4797 = _GEN_6085 == 10'h324 ? _GEN_4796 : _GEN_4795; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4798 = ~io_inputBit ? 1'h0 : _GEN_4797; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4799 = _GEN_6085 == 10'h325 ? _GEN_4798 : _GEN_4797; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4800 = io_inputBit | _GEN_4799; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4801 = _GEN_6085 == 10'h325 ? _GEN_4800 : _GEN_4799; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4802 = ~io_inputBit ? 1'h0 : _GEN_4801; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4803 = _GEN_6085 == 10'h326 ? _GEN_4802 : _GEN_4801; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4804 = io_inputBit | _GEN_4803; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4805 = _GEN_6085 == 10'h326 ? _GEN_4804 : _GEN_4803; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4806 = ~io_inputBit ? 1'h0 : _GEN_4805; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4807 = _GEN_6085 == 10'h327 ? _GEN_4806 : _GEN_4805; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4808 = io_inputBit | _GEN_4807; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4809 = _GEN_6085 == 10'h327 ? _GEN_4808 : _GEN_4807; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4810 = ~io_inputBit ? 1'h0 : _GEN_4809; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4811 = _GEN_6085 == 10'h328 ? _GEN_4810 : _GEN_4809; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4812 = io_inputBit | _GEN_4811; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4813 = _GEN_6085 == 10'h328 ? _GEN_4812 : _GEN_4811; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4814 = ~io_inputBit ? 1'h0 : _GEN_4813; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4815 = _GEN_6085 == 10'h329 ? _GEN_4814 : _GEN_4813; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4816 = io_inputBit | _GEN_4815; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4817 = _GEN_6085 == 10'h329 ? _GEN_4816 : _GEN_4815; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4818 = ~io_inputBit ? 1'h0 : _GEN_4817; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4819 = _GEN_6085 == 10'h32a ? _GEN_4818 : _GEN_4817; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4820 = io_inputBit | _GEN_4819; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4821 = _GEN_6085 == 10'h32a ? _GEN_4820 : _GEN_4819; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4822 = io_inputBit ? 1'h0 : _GEN_4269; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4823 = i == 8'h0 ? _GEN_4822 : _GEN_4269; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4824 = io_inputBit ? 1'h0 : _GEN_4823; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4825 = i == 8'h1 ? _GEN_4824 : _GEN_4823; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4826 = io_inputBit ? 1'h0 : _GEN_4825; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4827 = i == 8'h3 ? _GEN_4826 : _GEN_4825; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4828 = ~io_inputBit | _GEN_4827; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4829 = i == 8'h7 ? _GEN_4828 : _GEN_4827; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4830 = ~io_inputBit | _GEN_4829; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4831 = i == 8'h10 ? _GEN_4830 : _GEN_4829; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4832 = ~io_inputBit | _GEN_4831; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4833 = i == 8'h22 ? _GEN_4832 : _GEN_4831; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4834 = io_inputBit ? 1'h0 : _GEN_4833; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4835 = i == 8'h22 ? _GEN_4834 : _GEN_4833; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4836 = io_inputBit ? 1'h0 : _GEN_4301; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4837 = i == 8'h0 ? _GEN_4836 : _GEN_4301; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4838 = io_inputBit ? 1'h0 : _GEN_4837; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4839 = i == 8'h1 ? _GEN_4838 : _GEN_4837; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4840 = ~io_inputBit | _GEN_4839; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4841 = i == 8'h7 ? _GEN_4840 : _GEN_4839; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4842 = io_inputBit ? 1'h0 : _GEN_4841; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4843 = i == 8'h8 ? _GEN_4842 : _GEN_4841; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4844 = io_inputBit ? 1'h0 : _GEN_4843; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4845 = i == 8'h11 ? _GEN_4844 : _GEN_4843; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4846 = ~io_inputBit | _GEN_4845; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4847 = i == 8'h21 ? _GEN_4846 : _GEN_4845; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4848 = ~io_inputBit ? 1'h0 : _GEN_4847; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4849 = i == 8'h22 ? _GEN_4848 : _GEN_4847; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4850 = io_inputBit | _GEN_4849; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4851 = i == 8'h22 ? _GEN_4850 : _GEN_4849; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4852 = io_inputBit ? 1'h0 : _GEN_4851; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4853 = i == 8'h23 ? _GEN_4852 : _GEN_4851; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4854 = io_inputBit ? 1'h0 : _GEN_4853; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4855 = i == 8'h44 ? _GEN_4854 : _GEN_4853; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4856 = ~io_inputBit | _GEN_4855; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4857 = i == 8'h47 ? _GEN_4856 : _GEN_4855; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4858 = io_inputBit ? 1'h0 : _GEN_4857; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4859 = i == 8'h47 ? _GEN_4858 : _GEN_4857; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4860 = ~io_inputBit | _GEN_4859; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4861 = i == 8'h89 ? _GEN_4860 : _GEN_4859; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4862 = io_inputBit ? 1'h0 : _GEN_4861; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4863 = i == 8'h89 ? _GEN_4862 : _GEN_4861; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4864 = io_inputBit ? 1'h0 : _GEN_4345; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4865 = i == 8'h0 ? _GEN_4864 : _GEN_4345; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4866 = io_inputBit ? 1'h0 : _GEN_4865; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4867 = i == 8'h1 ? _GEN_4866 : _GEN_4865; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4868 = ~io_inputBit ? 1'h0 : _GEN_4867; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4869 = i == 8'h7 ? _GEN_4868 : _GEN_4867; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4870 = io_inputBit ? 1'h0 : _GEN_4869; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4871 = i == 8'h8 ? _GEN_4870 : _GEN_4869; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4872 = io_inputBit ? 1'h0 : _GEN_4871; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4873 = i == 8'h11 ? _GEN_4872 : _GEN_4871; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4874 = ~io_inputBit ? 1'h0 : _GEN_4873; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4875 = i == 8'h21 ? _GEN_4874 : _GEN_4873; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4876 = io_inputBit | _GEN_4875; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4877 = i == 8'h44 ? _GEN_4876 : _GEN_4875; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4878 = io_inputBit ? 1'h0 : _GEN_4877; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4879 = i == 8'h45 ? _GEN_4878 : _GEN_4877; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4880 = ~io_inputBit | _GEN_4879; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4881 = i == 8'h46 ? _GEN_4880 : _GEN_4879; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4882 = ~io_inputBit ? 1'h0 : _GEN_4881; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4883 = i == 8'h47 ? _GEN_4882 : _GEN_4881; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4884 = io_inputBit | _GEN_4883; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4885 = i == 8'h47 ? _GEN_4884 : _GEN_4883; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4886 = io_inputBit ? 1'h0 : _GEN_4885; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4887 = i == 8'h48 ? _GEN_4886 : _GEN_4885; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4888 = ~io_inputBit ? 1'h0 : _GEN_4887; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4889 = i == 8'h89 ? _GEN_4888 : _GEN_4887; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4890 = io_inputBit | _GEN_4889; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4891 = i == 8'h89 ? _GEN_4890 : _GEN_4889; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4892 = ~io_inputBit | _GEN_4891; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4893 = i == 8'h8b ? _GEN_4892 : _GEN_4891; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4894 = io_inputBit ? 1'h0 : _GEN_4893; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4895 = i == 8'h8b ? _GEN_4894 : _GEN_4893; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4896 = ~io_inputBit | _GEN_4895; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4897 = i == 8'h8e ? _GEN_4896 : _GEN_4895; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4898 = io_inputBit ? 1'h0 : _GEN_4897; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4899 = i == 8'h8e ? _GEN_4898 : _GEN_4897; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4900 = ~io_inputBit | _GEN_4899; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4901 = i == 8'h91 ? _GEN_4900 : _GEN_4899; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4902 = io_inputBit ? 1'h0 : _GEN_4901; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4903 = i == 8'h91 ? _GEN_4902 : _GEN_4901; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4904 = io_inputBit ? 1'h0 : _GEN_4413; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4905 = i == 8'h0 ? _GEN_4904 : _GEN_4413; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4906 = io_inputBit ? 1'h0 : _GEN_4905; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4907 = i == 8'h1 ? _GEN_4906 : _GEN_4905; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4908 = ~io_inputBit ? 1'h0 : _GEN_4907; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4909 = i == 8'h7 ? _GEN_4908 : _GEN_4907; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4910 = io_inputBit ? 1'h0 : _GEN_4909; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4911 = i == 8'h8 ? _GEN_4910 : _GEN_4909; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4912 = io_inputBit ? 1'h0 : _GEN_4911; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4913 = i == 8'h11 ? _GEN_4912 : _GEN_4911; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4914 = ~io_inputBit ? 1'h0 : _GEN_4913; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4915 = i == 8'h21 ? _GEN_4914 : _GEN_4913; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4916 = io_inputBit ? 1'h0 : _GEN_4915; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4917 = i == 8'h45 ? _GEN_4916 : _GEN_4915; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4918 = io_inputBit | _GEN_4917; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4919 = i == 8'h47 ? _GEN_4918 : _GEN_4917; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4920 = ~io_inputBit ? 1'h0 : _GEN_4919; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4921 = i == 8'h89 ? _GEN_4920 : _GEN_4919; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4922 = io_inputBit | _GEN_4921; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4923 = i == 8'h89 ? _GEN_4922 : _GEN_4921; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4924 = ~io_inputBit | _GEN_4923; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4925 = i == 8'h8a ? _GEN_4924 : _GEN_4923; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4926 = io_inputBit ? 1'h0 : _GEN_4925; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4927 = i == 8'h8a ? _GEN_4926 : _GEN_4925; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4928 = ~io_inputBit ? 1'h0 : _GEN_4927; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4929 = i == 8'h8b ? _GEN_4928 : _GEN_4927; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4930 = io_inputBit | _GEN_4929; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4931 = i == 8'h8b ? _GEN_4930 : _GEN_4929; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4932 = ~io_inputBit | _GEN_4931; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4933 = i == 8'h8d ? _GEN_4932 : _GEN_4931; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4934 = io_inputBit ? 1'h0 : _GEN_4933; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4935 = i == 8'h8d ? _GEN_4934 : _GEN_4933; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4936 = ~io_inputBit ? 1'h0 : _GEN_4935; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4937 = i == 8'h8e ? _GEN_4936 : _GEN_4935; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4938 = io_inputBit | _GEN_4937; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4939 = i == 8'h8e ? _GEN_4938 : _GEN_4937; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4940 = ~io_inputBit | _GEN_4939; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4941 = i == 8'h8f ? _GEN_4940 : _GEN_4939; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4942 = io_inputBit ? 1'h0 : _GEN_4941; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4943 = i == 8'h8f ? _GEN_4942 : _GEN_4941; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4944 = ~io_inputBit ? 1'h0 : _GEN_4943; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4945 = i == 8'h91 ? _GEN_4944 : _GEN_4943; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4946 = io_inputBit | _GEN_4945; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4947 = i == 8'h91 ? _GEN_4946 : _GEN_4945; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4948 = ~io_inputBit | _GEN_4947; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4949 = i == 8'h92 ? _GEN_4948 : _GEN_4947; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4950 = io_inputBit ? 1'h0 : _GEN_4949; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4951 = i == 8'h92 ? _GEN_4950 : _GEN_4949; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4952 = io_inputBit ? 1'h0 : _GEN_4481; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4953 = i == 8'h0 ? _GEN_4952 : _GEN_4481; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4954 = io_inputBit ? 1'h0 : _GEN_4953; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4955 = i == 8'h1 ? _GEN_4954 : _GEN_4953; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4956 = ~io_inputBit | _GEN_4955; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4957 = i == 8'h7 ? _GEN_4956 : _GEN_4955; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4958 = io_inputBit ? 1'h0 : _GEN_4957; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4959 = i == 8'h8 ? _GEN_4958 : _GEN_4957; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4960 = io_inputBit ? 1'h0 : _GEN_4959; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4961 = i == 8'h11 ? _GEN_4960 : _GEN_4959; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4962 = ~io_inputBit | _GEN_4961; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4963 = i == 8'h21 ? _GEN_4962 : _GEN_4961; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4964 = ~io_inputBit | _GEN_4963; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4965 = i == 8'h44 ? _GEN_4964 : _GEN_4963; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4966 = ~io_inputBit ? 1'h0 : _GEN_4965; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4967 = i == 8'h45 ? _GEN_4966 : _GEN_4965; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4968 = ~io_inputBit | _GEN_4967; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4969 = i == 8'h46 ? _GEN_4968 : _GEN_4967; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4970 = ~io_inputBit ? 1'h0 : _GEN_4969; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4971 = i == 8'h47 ? _GEN_4970 : _GEN_4969; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4972 = ~io_inputBit | _GEN_4971; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4973 = i == 8'h48 ? _GEN_4972 : _GEN_4971; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4974 = ~io_inputBit ? 1'h0 : _GEN_4973; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4975 = i == 8'h8a ? _GEN_4974 : _GEN_4973; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4976 = io_inputBit | _GEN_4975; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4977 = i == 8'h8a ? _GEN_4976 : _GEN_4975; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4978 = ~io_inputBit | _GEN_4977; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4979 = i == 8'h8c ? _GEN_4978 : _GEN_4977; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4980 = io_inputBit ? 1'h0 : _GEN_4979; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4981 = i == 8'h8c ? _GEN_4980 : _GEN_4979; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4982 = ~io_inputBit ? 1'h0 : _GEN_4981; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4983 = i == 8'h8e ? _GEN_4982 : _GEN_4981; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4984 = io_inputBit | _GEN_4983; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4985 = i == 8'h8e ? _GEN_4984 : _GEN_4983; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4986 = ~io_inputBit | _GEN_4985; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4987 = i == 8'h90 ? _GEN_4986 : _GEN_4985; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4988 = io_inputBit ? 1'h0 : _GEN_4987; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4989 = i == 8'h90 ? _GEN_4988 : _GEN_4987; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4990 = ~io_inputBit ? 1'h0 : _GEN_4989; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4991 = i == 8'h92 ? _GEN_4990 : _GEN_4989; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4992 = io_inputBit | _GEN_4991; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4993 = i == 8'h92 ? _GEN_4992 : _GEN_4991; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4994 = io_inputBit ? 1'h0 : _GEN_4601; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4995 = i == 8'h0 ? _GEN_4994 : _GEN_4601; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4996 = io_inputBit ? 1'h0 : _GEN_4995; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4997 = i == 8'h1 ? _GEN_4996 : _GEN_4995; // @[lut_mem_online.scala 235:34]
  wire  _GEN_4998 = ~io_inputBit ? 1'h0 : _GEN_4997; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_4999 = i == 8'h7 ? _GEN_4998 : _GEN_4997; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5000 = io_inputBit ? 1'h0 : _GEN_4999; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5001 = i == 8'h8 ? _GEN_5000 : _GEN_4999; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5002 = io_inputBit ? 1'h0 : _GEN_5001; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5003 = i == 8'h11 ? _GEN_5002 : _GEN_5001; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5004 = ~io_inputBit ? 1'h0 : _GEN_5003; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5005 = i == 8'h21 ? _GEN_5004 : _GEN_5003; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5006 = ~io_inputBit ? 1'h0 : _GEN_5005; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5007 = i == 8'h89 ? _GEN_5006 : _GEN_5005; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5008 = io_inputBit | _GEN_5007; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5009 = i == 8'h89 ? _GEN_5008 : _GEN_5007; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5010 = ~io_inputBit | _GEN_5009; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5011 = i == 8'h8a ? _GEN_5010 : _GEN_5009; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5012 = io_inputBit ? 1'h0 : _GEN_5011; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5013 = i == 8'h8a ? _GEN_5012 : _GEN_5011; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5014 = ~io_inputBit ? 1'h0 : _GEN_5013; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5015 = i == 8'h8b ? _GEN_5014 : _GEN_5013; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5016 = io_inputBit | _GEN_5015; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5017 = i == 8'h8b ? _GEN_5016 : _GEN_5015; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5018 = ~io_inputBit | _GEN_5017; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5019 = i == 8'h8c ? _GEN_5018 : _GEN_5017; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5020 = io_inputBit ? 1'h0 : _GEN_5019; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5021 = i == 8'h8c ? _GEN_5020 : _GEN_5019; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5022 = ~io_inputBit ? 1'h0 : _GEN_5021; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5023 = i == 8'h8d ? _GEN_5022 : _GEN_5021; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5024 = io_inputBit | _GEN_5023; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5025 = i == 8'h8d ? _GEN_5024 : _GEN_5023; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5026 = ~io_inputBit | _GEN_5025; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5027 = i == 8'h8e ? _GEN_5026 : _GEN_5025; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5028 = io_inputBit ? 1'h0 : _GEN_5027; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5029 = i == 8'h8e ? _GEN_5028 : _GEN_5027; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5030 = ~io_inputBit ? 1'h0 : _GEN_5029; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5031 = i == 8'h8f ? _GEN_5030 : _GEN_5029; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5032 = io_inputBit | _GEN_5031; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5033 = i == 8'h8f ? _GEN_5032 : _GEN_5031; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5034 = ~io_inputBit | _GEN_5033; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5035 = i == 8'h90 ? _GEN_5034 : _GEN_5033; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5036 = io_inputBit ? 1'h0 : _GEN_5035; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5037 = i == 8'h90 ? _GEN_5036 : _GEN_5035; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5038 = ~io_inputBit ? 1'h0 : _GEN_5037; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5039 = i == 8'h91 ? _GEN_5038 : _GEN_5037; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5040 = io_inputBit | _GEN_5039; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5041 = i == 8'h91 ? _GEN_5040 : _GEN_5039; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5042 = ~io_inputBit | _GEN_5041; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5043 = i == 8'h92 ? _GEN_5042 : _GEN_5041; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5044 = io_inputBit ? 1'h0 : _GEN_5043; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5045 = i == 8'h92 ? _GEN_5044 : _GEN_5043; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5046 = io_inputBit ? 1'h0 : _GEN_4821; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5047 = i == 8'h0 ? _GEN_5046 : _GEN_4821; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5048 = io_inputBit ? 1'h0 : _GEN_5047; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5049 = i == 8'h1 ? _GEN_5048 : _GEN_5047; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5050 = ~io_inputBit ? 1'h0 : _GEN_5049; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5051 = i == 8'h7 ? _GEN_5050 : _GEN_5049; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5052 = io_inputBit ? 1'h0 : _GEN_5051; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5053 = i == 8'h8 ? _GEN_5052 : _GEN_5051; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5054 = io_inputBit ? 1'h0 : _GEN_5053; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5055 = i == 8'h11 ? _GEN_5054 : _GEN_5053; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5056 = ~io_inputBit ? 1'h0 : _GEN_5055; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5057 = i == 8'h21 ? _GEN_5056 : _GEN_5055; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5058 = ~io_inputBit ? 1'h0 : _GEN_5057; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5059 = i == 8'h89 ? _GEN_5058 : _GEN_5057; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5060 = io_inputBit | _GEN_5059; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5061 = i == 8'h89 ? _GEN_5060 : _GEN_5059; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5062 = ~io_inputBit ? 1'h0 : _GEN_5061; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5063 = i == 8'h8a ? _GEN_5062 : _GEN_5061; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5064 = io_inputBit | _GEN_5063; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5065 = i == 8'h8a ? _GEN_5064 : _GEN_5063; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5066 = ~io_inputBit ? 1'h0 : _GEN_5065; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5067 = i == 8'h8b ? _GEN_5066 : _GEN_5065; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5068 = io_inputBit | _GEN_5067; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5069 = i == 8'h8b ? _GEN_5068 : _GEN_5067; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5070 = ~io_inputBit ? 1'h0 : _GEN_5069; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5071 = i == 8'h8c ? _GEN_5070 : _GEN_5069; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5072 = io_inputBit | _GEN_5071; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5073 = i == 8'h8c ? _GEN_5072 : _GEN_5071; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5074 = ~io_inputBit ? 1'h0 : _GEN_5073; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5075 = i == 8'h8d ? _GEN_5074 : _GEN_5073; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5076 = io_inputBit | _GEN_5075; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5077 = i == 8'h8d ? _GEN_5076 : _GEN_5075; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5078 = ~io_inputBit ? 1'h0 : _GEN_5077; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5079 = i == 8'h8e ? _GEN_5078 : _GEN_5077; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5080 = io_inputBit | _GEN_5079; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5081 = i == 8'h8e ? _GEN_5080 : _GEN_5079; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5082 = ~io_inputBit ? 1'h0 : _GEN_5081; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5083 = i == 8'h8f ? _GEN_5082 : _GEN_5081; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5084 = io_inputBit | _GEN_5083; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5085 = i == 8'h8f ? _GEN_5084 : _GEN_5083; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5086 = ~io_inputBit ? 1'h0 : _GEN_5085; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5087 = i == 8'h90 ? _GEN_5086 : _GEN_5085; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5088 = io_inputBit | _GEN_5087; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5089 = i == 8'h90 ? _GEN_5088 : _GEN_5087; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5090 = ~io_inputBit ? 1'h0 : _GEN_5089; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5091 = i == 8'h91 ? _GEN_5090 : _GEN_5089; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5092 = io_inputBit | _GEN_5091; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5093 = i == 8'h91 ? _GEN_5092 : _GEN_5091; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5094 = ~io_inputBit ? 1'h0 : _GEN_5093; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5095 = i == 8'h92 ? _GEN_5094 : _GEN_5093; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5096 = io_inputBit | _GEN_5095; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5097 = i == 8'h92 ? _GEN_5096 : _GEN_5095; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5098 = io_inputBit ? 1'h0 : _GEN_4835; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5099 = i == 8'h0 ? _GEN_5098 : _GEN_4835; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5100 = ~io_inputBit ? 1'h0 : _GEN_5099; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5101 = i == 8'h3 ? _GEN_5100 : _GEN_5099; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5102 = io_inputBit ? 1'h0 : _GEN_5101; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5103 = i == 8'h4 ? _GEN_5102 : _GEN_5101; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5104 = io_inputBit | _GEN_5103; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5105 = i == 8'h8 ? _GEN_5104 : _GEN_5103; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5106 = io_inputBit ? 1'h0 : _GEN_5105; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5107 = i == 8'h9 ? _GEN_5106 : _GEN_5105; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5108 = io_inputBit | _GEN_5107; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5109 = i == 8'h11 ? _GEN_5108 : _GEN_5107; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5110 = io_inputBit ? 1'h0 : _GEN_5109; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5111 = i == 8'h13 ? _GEN_5110 : _GEN_5109; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5112 = io_inputBit | _GEN_5111; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5113 = i == 8'h23 ? _GEN_5112 : _GEN_5111; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5114 = ~io_inputBit | _GEN_5113; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5115 = i == 8'h27 ? _GEN_5114 : _GEN_5113; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5116 = io_inputBit ? 1'h0 : _GEN_5115; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5117 = i == 8'h27 ? _GEN_5116 : _GEN_5115; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5118 = io_inputBit | _GEN_5117; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5119 = i == 8'h47 ? _GEN_5118 : _GEN_5117; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5120 = ~io_inputBit ? 1'h0 : _GEN_5119; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5121 = i == 8'h8f ? _GEN_5120 : _GEN_5119; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5122 = io_inputBit | _GEN_5121; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5123 = i == 8'h8f ? _GEN_5122 : _GEN_5121; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5124 = io_inputBit ? 1'h0 : _GEN_4863; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5125 = i == 8'h0 ? _GEN_5124 : _GEN_4863; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5126 = io_inputBit ? 1'h0 : _GEN_5125; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5127 = i == 8'h4 ? _GEN_5126 : _GEN_5125; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5128 = ~io_inputBit ? 1'h0 : _GEN_5127; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5129 = i == 8'h7 ? _GEN_5128 : _GEN_5127; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5130 = io_inputBit ? 1'h0 : _GEN_5129; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5131 = i == 8'h9 ? _GEN_5130 : _GEN_5129; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5132 = ~io_inputBit ? 1'h0 : _GEN_5131; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5133 = i == 8'h10 ? _GEN_5132 : _GEN_5131; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5134 = io_inputBit | _GEN_5133; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5135 = i == 8'h11 ? _GEN_5134 : _GEN_5133; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5136 = ~io_inputBit | _GEN_5135; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5137 = i == 8'h12 ? _GEN_5136 : _GEN_5135; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5138 = io_inputBit | _GEN_5137; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5139 = i == 8'h22 ? _GEN_5138 : _GEN_5137; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5140 = io_inputBit ? 1'h0 : _GEN_5139; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5141 = i == 8'h23 ? _GEN_5140 : _GEN_5139; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5142 = ~io_inputBit | _GEN_5141; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5143 = i == 8'h26 ? _GEN_5142 : _GEN_5141; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5144 = ~io_inputBit ? 1'h0 : _GEN_5143; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5145 = i == 8'h27 ? _GEN_5144 : _GEN_5143; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5146 = io_inputBit | _GEN_5145; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5147 = i == 8'h27 ? _GEN_5146 : _GEN_5145; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5148 = io_inputBit ? 1'h0 : _GEN_5147; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5149 = i == 8'h28 ? _GEN_5148 : _GEN_5147; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5150 = ~io_inputBit ? 1'h0 : _GEN_5149; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5151 = i == 8'h45 ? _GEN_5150 : _GEN_5149; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5152 = io_inputBit ? 1'h0 : _GEN_5151; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5153 = i == 8'h47 ? _GEN_5152 : _GEN_5151; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5154 = io_inputBit ? 1'h0 : _GEN_5153; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5155 = i == 8'h4e ? _GEN_5154 : _GEN_5153; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5156 = ~io_inputBit | _GEN_5155; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5157 = i == 8'h51 ? _GEN_5156 : _GEN_5155; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5158 = io_inputBit ? 1'h0 : _GEN_5157; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5159 = i == 8'h51 ? _GEN_5158 : _GEN_5157; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5160 = ~io_inputBit ? 1'h0 : _GEN_5159; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5161 = i == 8'h8c ? _GEN_5160 : _GEN_5159; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5162 = io_inputBit | _GEN_5161; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5163 = i == 8'h8c ? _GEN_5162 : _GEN_5161; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5164 = ~io_inputBit | _GEN_5163; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5165 = i == 8'h8f ? _GEN_5164 : _GEN_5163; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5166 = io_inputBit ? 1'h0 : _GEN_5165; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5167 = i == 8'h8f ? _GEN_5166 : _GEN_5165; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5168 = ~io_inputBit | _GEN_5167; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5169 = i == 8'h9d ? _GEN_5168 : _GEN_5167; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5170 = io_inputBit ? 1'h0 : _GEN_5169; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5171 = i == 8'h9d ? _GEN_5170 : _GEN_5169; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5172 = io_inputBit ? 1'h0 : _GEN_4903; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5173 = i == 8'h0 ? _GEN_5172 : _GEN_4903; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5174 = io_inputBit ? 1'h0 : _GEN_5173; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5175 = i == 8'h4 ? _GEN_5174 : _GEN_5173; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5176 = ~io_inputBit ? 1'h0 : _GEN_5175; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5177 = i == 8'h7 ? _GEN_5176 : _GEN_5175; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5178 = io_inputBit ? 1'h0 : _GEN_5177; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5179 = i == 8'h9 ? _GEN_5178 : _GEN_5177; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5180 = ~io_inputBit ? 1'h0 : _GEN_5179; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5181 = i == 8'h10 ? _GEN_5180 : _GEN_5179; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5182 = io_inputBit ? 1'h0 : _GEN_5181; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5183 = i == 8'h11 ? _GEN_5182 : _GEN_5181; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5184 = ~io_inputBit ? 1'h0 : _GEN_5183; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5185 = i == 8'h12 ? _GEN_5184 : _GEN_5183; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5186 = io_inputBit | _GEN_5185; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5187 = i == 8'h23 ? _GEN_5186 : _GEN_5185; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5188 = ~io_inputBit ? 1'h0 : _GEN_5187; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5189 = i == 8'h26 ? _GEN_5188 : _GEN_5187; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5190 = ~io_inputBit | _GEN_5189; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5191 = i == 8'h45 ? _GEN_5190 : _GEN_5189; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5192 = ~io_inputBit ? 1'h0 : _GEN_5191; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5193 = i == 8'h46 ? _GEN_5192 : _GEN_5191; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5194 = io_inputBit | _GEN_5193; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5195 = i == 8'h46 ? _GEN_5194 : _GEN_5193; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5196 = io_inputBit ? 1'h0 : _GEN_5195; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5197 = i == 8'h47 ? _GEN_5196 : _GEN_5195; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5198 = io_inputBit | _GEN_5197; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5199 = i == 8'h4e ? _GEN_5198 : _GEN_5197; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5200 = io_inputBit ? 1'h0 : _GEN_5199; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5201 = i == 8'h4f ? _GEN_5200 : _GEN_5199; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5202 = ~io_inputBit | _GEN_5201; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5203 = i == 8'h50 ? _GEN_5202 : _GEN_5201; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5204 = ~io_inputBit ? 1'h0 : _GEN_5203; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5205 = i == 8'h51 ? _GEN_5204 : _GEN_5203; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5206 = io_inputBit | _GEN_5205; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5207 = i == 8'h51 ? _GEN_5206 : _GEN_5205; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5208 = io_inputBit ? 1'h0 : _GEN_5207; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5209 = i == 8'h52 ? _GEN_5208 : _GEN_5207; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5210 = ~io_inputBit | _GEN_5209; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5211 = i == 8'h8c ? _GEN_5210 : _GEN_5209; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5212 = io_inputBit ? 1'h0 : _GEN_5211; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5213 = i == 8'h8c ? _GEN_5212 : _GEN_5211; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5214 = ~io_inputBit | _GEN_5213; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5215 = i == 8'h8f ? _GEN_5214 : _GEN_5213; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5216 = io_inputBit ? 1'h0 : _GEN_5215; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5217 = i == 8'h8f ? _GEN_5216 : _GEN_5215; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5218 = ~io_inputBit ? 1'h0 : _GEN_5217; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5219 = i == 8'h9d ? _GEN_5218 : _GEN_5217; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5220 = io_inputBit | _GEN_5219; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5221 = i == 8'h9d ? _GEN_5220 : _GEN_5219; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5222 = ~io_inputBit | _GEN_5221; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5223 = i == 8'h9f ? _GEN_5222 : _GEN_5221; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5224 = io_inputBit ? 1'h0 : _GEN_5223; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5225 = i == 8'h9f ? _GEN_5224 : _GEN_5223; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5226 = ~io_inputBit | _GEN_5225; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5227 = i == 8'ha2 ? _GEN_5226 : _GEN_5225; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5228 = io_inputBit ? 1'h0 : _GEN_5227; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5229 = i == 8'ha2 ? _GEN_5228 : _GEN_5227; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5230 = ~io_inputBit | _GEN_5229; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5231 = i == 8'ha5 ? _GEN_5230 : _GEN_5229; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5232 = io_inputBit ? 1'h0 : _GEN_5231; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5233 = i == 8'ha5 ? _GEN_5232 : _GEN_5231; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5234 = io_inputBit ? 1'h0 : _GEN_4951; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5235 = i == 8'h0 ? _GEN_5234 : _GEN_4951; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5236 = io_inputBit ? 1'h0 : _GEN_5235; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5237 = i == 8'h4 ? _GEN_5236 : _GEN_5235; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5238 = ~io_inputBit ? 1'h0 : _GEN_5237; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5239 = i == 8'h7 ? _GEN_5238 : _GEN_5237; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5240 = io_inputBit ? 1'h0 : _GEN_5239; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5241 = i == 8'h9 ? _GEN_5240 : _GEN_5239; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5242 = io_inputBit ? 1'h0 : _GEN_5241; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5243 = i == 8'h11 ? _GEN_5242 : _GEN_5241; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5244 = ~io_inputBit ? 1'h0 : _GEN_5243; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5245 = i == 8'h12 ? _GEN_5244 : _GEN_5243; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5246 = ~io_inputBit ? 1'h0 : _GEN_5245; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5247 = i == 8'h21 ? _GEN_5246 : _GEN_5245; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5248 = ~io_inputBit ? 1'h0 : _GEN_5247; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5249 = i == 8'h26 ? _GEN_5248 : _GEN_5247; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5250 = ~io_inputBit ? 1'h0 : _GEN_5249; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5251 = i == 8'h44 ? _GEN_5250 : _GEN_5249; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5252 = io_inputBit | _GEN_5251; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5253 = i == 8'h44 ? _GEN_5252 : _GEN_5251; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5254 = ~io_inputBit | _GEN_5253; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5255 = i == 8'h46 ? _GEN_5254 : _GEN_5253; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5256 = io_inputBit ? 1'h0 : _GEN_5255; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5257 = i == 8'h46 ? _GEN_5256 : _GEN_5255; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5258 = ~io_inputBit ? 1'h0 : _GEN_5257; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5259 = i == 8'h48 ? _GEN_5258 : _GEN_5257; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5260 = io_inputBit | _GEN_5259; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5261 = i == 8'h48 ? _GEN_5260 : _GEN_5259; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5262 = io_inputBit ? 1'h0 : _GEN_5261; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5263 = i == 8'h4f ? _GEN_5262 : _GEN_5261; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5264 = io_inputBit | _GEN_5263; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5265 = i == 8'h51 ? _GEN_5264 : _GEN_5263; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5266 = ~io_inputBit ? 1'h0 : _GEN_5265; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5267 = i == 8'h8b ? _GEN_5266 : _GEN_5265; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5268 = io_inputBit | _GEN_5267; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5269 = i == 8'h8b ? _GEN_5268 : _GEN_5267; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5270 = ~io_inputBit | _GEN_5269; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5271 = i == 8'h8c ? _GEN_5270 : _GEN_5269; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5272 = io_inputBit ? 1'h0 : _GEN_5271; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5273 = i == 8'h8c ? _GEN_5272 : _GEN_5271; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5274 = ~io_inputBit | _GEN_5273; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5275 = i == 8'h8f ? _GEN_5274 : _GEN_5273; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5276 = io_inputBit ? 1'h0 : _GEN_5275; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5277 = i == 8'h8f ? _GEN_5276 : _GEN_5275; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5278 = ~io_inputBit ? 1'h0 : _GEN_5277; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5279 = i == 8'h90 ? _GEN_5278 : _GEN_5277; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5280 = io_inputBit | _GEN_5279; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5281 = i == 8'h90 ? _GEN_5280 : _GEN_5279; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5282 = ~io_inputBit ? 1'h0 : _GEN_5281; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5283 = i == 8'h9d ? _GEN_5282 : _GEN_5281; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5284 = io_inputBit | _GEN_5283; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5285 = i == 8'h9d ? _GEN_5284 : _GEN_5283; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5286 = ~io_inputBit | _GEN_5285; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5287 = i == 8'h9e ? _GEN_5286 : _GEN_5285; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5288 = io_inputBit ? 1'h0 : _GEN_5287; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5289 = i == 8'h9e ? _GEN_5288 : _GEN_5287; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5290 = ~io_inputBit ? 1'h0 : _GEN_5289; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5291 = i == 8'h9f ? _GEN_5290 : _GEN_5289; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5292 = io_inputBit | _GEN_5291; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5293 = i == 8'h9f ? _GEN_5292 : _GEN_5291; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5294 = ~io_inputBit | _GEN_5293; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5295 = i == 8'ha1 ? _GEN_5294 : _GEN_5293; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5296 = io_inputBit ? 1'h0 : _GEN_5295; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5297 = i == 8'ha1 ? _GEN_5296 : _GEN_5295; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5298 = ~io_inputBit ? 1'h0 : _GEN_5297; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5299 = i == 8'ha2 ? _GEN_5298 : _GEN_5297; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5300 = io_inputBit | _GEN_5299; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5301 = i == 8'ha2 ? _GEN_5300 : _GEN_5299; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5302 = ~io_inputBit | _GEN_5301; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5303 = i == 8'ha3 ? _GEN_5302 : _GEN_5301; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5304 = io_inputBit ? 1'h0 : _GEN_5303; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5305 = i == 8'ha3 ? _GEN_5304 : _GEN_5303; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5306 = ~io_inputBit ? 1'h0 : _GEN_5305; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5307 = i == 8'ha5 ? _GEN_5306 : _GEN_5305; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5308 = io_inputBit | _GEN_5307; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5309 = i == 8'ha5 ? _GEN_5308 : _GEN_5307; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5310 = ~io_inputBit | _GEN_5309; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5311 = i == 8'ha6 ? _GEN_5310 : _GEN_5309; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5312 = io_inputBit ? 1'h0 : _GEN_5311; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5313 = i == 8'ha6 ? _GEN_5312 : _GEN_5311; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5314 = io_inputBit ? 1'h0 : _GEN_4993; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5315 = i == 8'h0 ? _GEN_5314 : _GEN_4993; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5316 = io_inputBit ? 1'h0 : _GEN_5315; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5317 = i == 8'h4 ? _GEN_5316 : _GEN_5315; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5318 = ~io_inputBit ? 1'h0 : _GEN_5317; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5319 = i == 8'h7 ? _GEN_5318 : _GEN_5317; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5320 = io_inputBit ? 1'h0 : _GEN_5319; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5321 = i == 8'h9 ? _GEN_5320 : _GEN_5319; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5322 = io_inputBit | _GEN_5321; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5323 = i == 8'h11 ? _GEN_5322 : _GEN_5321; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5324 = ~io_inputBit | _GEN_5323; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5325 = i == 8'h12 ? _GEN_5324 : _GEN_5323; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5326 = ~io_inputBit ? 1'h0 : _GEN_5325; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5327 = i == 8'h21 ? _GEN_5326 : _GEN_5325; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5328 = ~io_inputBit | _GEN_5327; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5329 = i == 8'h26 ? _GEN_5328 : _GEN_5327; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5330 = ~io_inputBit | _GEN_5329; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5331 = i == 8'h4e ? _GEN_5330 : _GEN_5329; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5332 = ~io_inputBit ? 1'h0 : _GEN_5331; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5333 = i == 8'h4f ? _GEN_5332 : _GEN_5331; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5334 = ~io_inputBit | _GEN_5333; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5335 = i == 8'h50 ? _GEN_5334 : _GEN_5333; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5336 = ~io_inputBit ? 1'h0 : _GEN_5335; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5337 = i == 8'h51 ? _GEN_5336 : _GEN_5335; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5338 = ~io_inputBit | _GEN_5337; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5339 = i == 8'h52 ? _GEN_5338 : _GEN_5337; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5340 = ~io_inputBit ? 1'h0 : _GEN_5339; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5341 = i == 8'h89 ? _GEN_5340 : _GEN_5339; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5342 = io_inputBit | _GEN_5341; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5343 = i == 8'h89 ? _GEN_5342 : _GEN_5341; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5344 = ~io_inputBit ? 1'h0 : _GEN_5343; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5345 = i == 8'h8a ? _GEN_5344 : _GEN_5343; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5346 = io_inputBit | _GEN_5345; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5347 = i == 8'h8a ? _GEN_5346 : _GEN_5345; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5348 = ~io_inputBit | _GEN_5347; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5349 = i == 8'h8b ? _GEN_5348 : _GEN_5347; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5350 = io_inputBit ? 1'h0 : _GEN_5349; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5351 = i == 8'h8b ? _GEN_5350 : _GEN_5349; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5352 = ~io_inputBit | _GEN_5351; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5353 = i == 8'h8c ? _GEN_5352 : _GEN_5351; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5354 = io_inputBit ? 1'h0 : _GEN_5353; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5355 = i == 8'h8c ? _GEN_5354 : _GEN_5353; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5356 = ~io_inputBit ? 1'h0 : _GEN_5355; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5357 = i == 8'h8d ? _GEN_5356 : _GEN_5355; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5358 = io_inputBit | _GEN_5357; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5359 = i == 8'h8d ? _GEN_5358 : _GEN_5357; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5360 = ~io_inputBit ? 1'h0 : _GEN_5359; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5361 = i == 8'h8e ? _GEN_5360 : _GEN_5359; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5362 = io_inputBit | _GEN_5361; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5363 = i == 8'h8e ? _GEN_5362 : _GEN_5361; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5364 = ~io_inputBit | _GEN_5363; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5365 = i == 8'h8f ? _GEN_5364 : _GEN_5363; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5366 = io_inputBit ? 1'h0 : _GEN_5365; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5367 = i == 8'h8f ? _GEN_5366 : _GEN_5365; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5368 = ~io_inputBit | _GEN_5367; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5369 = i == 8'h90 ? _GEN_5368 : _GEN_5367; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5370 = io_inputBit ? 1'h0 : _GEN_5369; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5371 = i == 8'h90 ? _GEN_5370 : _GEN_5369; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5372 = ~io_inputBit ? 1'h0 : _GEN_5371; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5373 = i == 8'h91 ? _GEN_5372 : _GEN_5371; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5374 = io_inputBit | _GEN_5373; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5375 = i == 8'h91 ? _GEN_5374 : _GEN_5373; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5376 = ~io_inputBit ? 1'h0 : _GEN_5375; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5377 = i == 8'h92 ? _GEN_5376 : _GEN_5375; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5378 = io_inputBit | _GEN_5377; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5379 = i == 8'h92 ? _GEN_5378 : _GEN_5377; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5380 = ~io_inputBit ? 1'h0 : _GEN_5379; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5381 = i == 8'h9e ? _GEN_5380 : _GEN_5379; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5382 = io_inputBit | _GEN_5381; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5383 = i == 8'h9e ? _GEN_5382 : _GEN_5381; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5384 = ~io_inputBit | _GEN_5383; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5385 = i == 8'ha0 ? _GEN_5384 : _GEN_5383; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5386 = io_inputBit ? 1'h0 : _GEN_5385; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5387 = i == 8'ha0 ? _GEN_5386 : _GEN_5385; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5388 = ~io_inputBit ? 1'h0 : _GEN_5387; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5389 = i == 8'ha2 ? _GEN_5388 : _GEN_5387; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5390 = io_inputBit | _GEN_5389; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5391 = i == 8'ha2 ? _GEN_5390 : _GEN_5389; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5392 = ~io_inputBit | _GEN_5391; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5393 = i == 8'ha4 ? _GEN_5392 : _GEN_5391; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5394 = io_inputBit ? 1'h0 : _GEN_5393; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5395 = i == 8'ha4 ? _GEN_5394 : _GEN_5393; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5396 = ~io_inputBit ? 1'h0 : _GEN_5395; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5397 = i == 8'ha6 ? _GEN_5396 : _GEN_5395; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5398 = io_inputBit | _GEN_5397; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5399 = i == 8'ha6 ? _GEN_5398 : _GEN_5397; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5400 = io_inputBit ? 1'h0 : _GEN_5045; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5401 = i == 8'h0 ? _GEN_5400 : _GEN_5045; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5402 = io_inputBit ? 1'h0 : _GEN_5401; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5403 = i == 8'h4 ? _GEN_5402 : _GEN_5401; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5404 = ~io_inputBit ? 1'h0 : _GEN_5403; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5405 = i == 8'h7 ? _GEN_5404 : _GEN_5403; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5406 = io_inputBit ? 1'h0 : _GEN_5405; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5407 = i == 8'h9 ? _GEN_5406 : _GEN_5405; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5408 = io_inputBit ? 1'h0 : _GEN_5407; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5409 = i == 8'h11 ? _GEN_5408 : _GEN_5407; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5410 = ~io_inputBit ? 1'h0 : _GEN_5409; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5411 = i == 8'h12 ? _GEN_5410 : _GEN_5409; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5412 = ~io_inputBit ? 1'h0 : _GEN_5411; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5413 = i == 8'h21 ? _GEN_5412 : _GEN_5411; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5414 = ~io_inputBit ? 1'h0 : _GEN_5413; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5415 = i == 8'h26 ? _GEN_5414 : _GEN_5413; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5416 = ~io_inputBit ? 1'h0 : _GEN_5415; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5417 = i == 8'h44 ? _GEN_5416 : _GEN_5415; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5418 = io_inputBit | _GEN_5417; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5419 = i == 8'h44 ? _GEN_5418 : _GEN_5417; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5420 = ~io_inputBit ? 1'h0 : _GEN_5419; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5421 = i == 8'h45 ? _GEN_5420 : _GEN_5419; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5422 = io_inputBit | _GEN_5421; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5423 = i == 8'h45 ? _GEN_5422 : _GEN_5421; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5424 = ~io_inputBit ? 1'h0 : _GEN_5423; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5425 = i == 8'h46 ? _GEN_5424 : _GEN_5423; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5426 = io_inputBit | _GEN_5425; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5427 = i == 8'h46 ? _GEN_5426 : _GEN_5425; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5428 = ~io_inputBit ? 1'h0 : _GEN_5427; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5429 = i == 8'h47 ? _GEN_5428 : _GEN_5427; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5430 = io_inputBit | _GEN_5429; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5431 = i == 8'h47 ? _GEN_5430 : _GEN_5429; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5432 = ~io_inputBit ? 1'h0 : _GEN_5431; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5433 = i == 8'h48 ? _GEN_5432 : _GEN_5431; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5434 = io_inputBit | _GEN_5433; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5435 = i == 8'h48 ? _GEN_5434 : _GEN_5433; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5436 = ~io_inputBit ? 1'h0 : _GEN_5435; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5437 = i == 8'h9d ? _GEN_5436 : _GEN_5435; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5438 = io_inputBit | _GEN_5437; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5439 = i == 8'h9d ? _GEN_5438 : _GEN_5437; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5440 = ~io_inputBit | _GEN_5439; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5441 = i == 8'h9e ? _GEN_5440 : _GEN_5439; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5442 = io_inputBit ? 1'h0 : _GEN_5441; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5443 = i == 8'h9e ? _GEN_5442 : _GEN_5441; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5444 = ~io_inputBit ? 1'h0 : _GEN_5443; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5445 = i == 8'h9f ? _GEN_5444 : _GEN_5443; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5446 = io_inputBit | _GEN_5445; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5447 = i == 8'h9f ? _GEN_5446 : _GEN_5445; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5448 = ~io_inputBit | _GEN_5447; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5449 = i == 8'ha0 ? _GEN_5448 : _GEN_5447; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5450 = io_inputBit ? 1'h0 : _GEN_5449; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5451 = i == 8'ha0 ? _GEN_5450 : _GEN_5449; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5452 = ~io_inputBit ? 1'h0 : _GEN_5451; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5453 = i == 8'ha1 ? _GEN_5452 : _GEN_5451; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5454 = io_inputBit | _GEN_5453; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5455 = i == 8'ha1 ? _GEN_5454 : _GEN_5453; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5456 = ~io_inputBit | _GEN_5455; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5457 = i == 8'ha2 ? _GEN_5456 : _GEN_5455; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5458 = io_inputBit ? 1'h0 : _GEN_5457; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5459 = i == 8'ha2 ? _GEN_5458 : _GEN_5457; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5460 = ~io_inputBit ? 1'h0 : _GEN_5459; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5461 = i == 8'ha3 ? _GEN_5460 : _GEN_5459; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5462 = io_inputBit | _GEN_5461; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5463 = i == 8'ha3 ? _GEN_5462 : _GEN_5461; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5464 = ~io_inputBit | _GEN_5463; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5465 = i == 8'ha4 ? _GEN_5464 : _GEN_5463; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5466 = io_inputBit ? 1'h0 : _GEN_5465; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5467 = i == 8'ha4 ? _GEN_5466 : _GEN_5465; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5468 = ~io_inputBit ? 1'h0 : _GEN_5467; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5469 = i == 8'ha5 ? _GEN_5468 : _GEN_5467; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5470 = io_inputBit | _GEN_5469; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5471 = i == 8'ha5 ? _GEN_5470 : _GEN_5469; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5472 = ~io_inputBit | _GEN_5471; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5473 = i == 8'ha6 ? _GEN_5472 : _GEN_5471; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5474 = io_inputBit ? 1'h0 : _GEN_5473; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5475 = i == 8'ha6 ? _GEN_5474 : _GEN_5473; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5476 = io_inputBit ? 1'h0 : _GEN_5097; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5477 = i == 8'h0 ? _GEN_5476 : _GEN_5097; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5478 = io_inputBit ? 1'h0 : _GEN_5477; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5479 = i == 8'h4 ? _GEN_5478 : _GEN_5477; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5480 = ~io_inputBit ? 1'h0 : _GEN_5479; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5481 = i == 8'h7 ? _GEN_5480 : _GEN_5479; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5482 = io_inputBit ? 1'h0 : _GEN_5481; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5483 = i == 8'h9 ? _GEN_5482 : _GEN_5481; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5484 = io_inputBit ? 1'h0 : _GEN_5483; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5485 = i == 8'h11 ? _GEN_5484 : _GEN_5483; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5486 = ~io_inputBit ? 1'h0 : _GEN_5485; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5487 = i == 8'h12 ? _GEN_5486 : _GEN_5485; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5488 = ~io_inputBit ? 1'h0 : _GEN_5487; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5489 = i == 8'h21 ? _GEN_5488 : _GEN_5487; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5490 = ~io_inputBit ? 1'h0 : _GEN_5489; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5491 = i == 8'h26 ? _GEN_5490 : _GEN_5489; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5492 = ~io_inputBit ? 1'h0 : _GEN_5491; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5493 = i == 8'h89 ? _GEN_5492 : _GEN_5491; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5494 = io_inputBit | _GEN_5493; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5495 = i == 8'h89 ? _GEN_5494 : _GEN_5493; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5496 = ~io_inputBit ? 1'h0 : _GEN_5495; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5497 = i == 8'h8a ? _GEN_5496 : _GEN_5495; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5498 = io_inputBit | _GEN_5497; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5499 = i == 8'h8a ? _GEN_5498 : _GEN_5497; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5500 = ~io_inputBit ? 1'h0 : _GEN_5499; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5501 = i == 8'h8b ? _GEN_5500 : _GEN_5499; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5502 = io_inputBit | _GEN_5501; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5503 = i == 8'h8b ? _GEN_5502 : _GEN_5501; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5504 = ~io_inputBit ? 1'h0 : _GEN_5503; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5505 = i == 8'h8c ? _GEN_5504 : _GEN_5503; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5506 = io_inputBit | _GEN_5505; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5507 = i == 8'h8c ? _GEN_5506 : _GEN_5505; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5508 = ~io_inputBit ? 1'h0 : _GEN_5507; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5509 = i == 8'h8d ? _GEN_5508 : _GEN_5507; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5510 = io_inputBit | _GEN_5509; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5511 = i == 8'h8d ? _GEN_5510 : _GEN_5509; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5512 = ~io_inputBit ? 1'h0 : _GEN_5511; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5513 = i == 8'h8e ? _GEN_5512 : _GEN_5511; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5514 = io_inputBit | _GEN_5513; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5515 = i == 8'h8e ? _GEN_5514 : _GEN_5513; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5516 = ~io_inputBit ? 1'h0 : _GEN_5515; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5517 = i == 8'h8f ? _GEN_5516 : _GEN_5515; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5518 = io_inputBit | _GEN_5517; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5519 = i == 8'h8f ? _GEN_5518 : _GEN_5517; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5520 = ~io_inputBit ? 1'h0 : _GEN_5519; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5521 = i == 8'h90 ? _GEN_5520 : _GEN_5519; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5522 = io_inputBit | _GEN_5521; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5523 = i == 8'h90 ? _GEN_5522 : _GEN_5521; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5524 = ~io_inputBit ? 1'h0 : _GEN_5523; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5525 = i == 8'h91 ? _GEN_5524 : _GEN_5523; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5526 = io_inputBit | _GEN_5525; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5527 = i == 8'h91 ? _GEN_5526 : _GEN_5525; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5528 = ~io_inputBit ? 1'h0 : _GEN_5527; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5529 = i == 8'h92 ? _GEN_5528 : _GEN_5527; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5530 = io_inputBit | _GEN_5529; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5531 = i == 8'h92 ? _GEN_5530 : _GEN_5529; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5532 = ~io_inputBit ? 1'h0 : _GEN_5531; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5533 = i == 8'h9d ? _GEN_5532 : _GEN_5531; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5534 = io_inputBit | _GEN_5533; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5535 = i == 8'h9d ? _GEN_5534 : _GEN_5533; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5536 = ~io_inputBit ? 1'h0 : _GEN_5535; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5537 = i == 8'h9e ? _GEN_5536 : _GEN_5535; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5538 = io_inputBit | _GEN_5537; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5539 = i == 8'h9e ? _GEN_5538 : _GEN_5537; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5540 = ~io_inputBit ? 1'h0 : _GEN_5539; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5541 = i == 8'h9f ? _GEN_5540 : _GEN_5539; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5542 = io_inputBit | _GEN_5541; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5543 = i == 8'h9f ? _GEN_5542 : _GEN_5541; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5544 = ~io_inputBit ? 1'h0 : _GEN_5543; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5545 = i == 8'ha0 ? _GEN_5544 : _GEN_5543; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5546 = io_inputBit | _GEN_5545; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5547 = i == 8'ha0 ? _GEN_5546 : _GEN_5545; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5548 = ~io_inputBit ? 1'h0 : _GEN_5547; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5549 = i == 8'ha1 ? _GEN_5548 : _GEN_5547; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5550 = io_inputBit | _GEN_5549; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5551 = i == 8'ha1 ? _GEN_5550 : _GEN_5549; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5552 = ~io_inputBit ? 1'h0 : _GEN_5551; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5553 = i == 8'ha2 ? _GEN_5552 : _GEN_5551; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5554 = io_inputBit | _GEN_5553; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5555 = i == 8'ha2 ? _GEN_5554 : _GEN_5553; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5556 = ~io_inputBit ? 1'h0 : _GEN_5555; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5557 = i == 8'ha3 ? _GEN_5556 : _GEN_5555; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5558 = io_inputBit | _GEN_5557; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5559 = i == 8'ha3 ? _GEN_5558 : _GEN_5557; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5560 = ~io_inputBit ? 1'h0 : _GEN_5559; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5561 = i == 8'ha4 ? _GEN_5560 : _GEN_5559; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5562 = io_inputBit | _GEN_5561; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5563 = i == 8'ha4 ? _GEN_5562 : _GEN_5561; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5564 = ~io_inputBit ? 1'h0 : _GEN_5563; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5565 = i == 8'ha5 ? _GEN_5564 : _GEN_5563; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5566 = io_inputBit | _GEN_5565; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5567 = i == 8'ha5 ? _GEN_5566 : _GEN_5565; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5568 = ~io_inputBit ? 1'h0 : _GEN_5567; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5569 = i == 8'ha6 ? _GEN_5568 : _GEN_5567; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5570 = io_inputBit | _GEN_5569; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5571 = i == 8'ha6 ? _GEN_5570 : _GEN_5569; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5572 = io_inputBit ? 1'h0 : _GEN_5123; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5573 = i == 8'h0 ? _GEN_5572 : _GEN_5123; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5574 = ~io_inputBit ? 1'h0 : _GEN_5573; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5575 = i == 8'h1 ? _GEN_5574 : _GEN_5573; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5576 = io_inputBit | _GEN_5575; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5577 = i == 8'h9 ? _GEN_5576 : _GEN_5575; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5578 = io_inputBit ? 1'h0 : _GEN_5577; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5579 = i == 8'ha ? _GEN_5578 : _GEN_5577; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5580 = ~io_inputBit ? 1'h0 : _GEN_5579; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5581 = i == 8'h13 ? _GEN_5580 : _GEN_5579; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5582 = ~io_inputBit | _GEN_5581; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5583 = i == 8'h15 ? _GEN_5582 : _GEN_5581; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5584 = io_inputBit | _GEN_5583; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5585 = i == 8'h28 ? _GEN_5584 : _GEN_5583; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5586 = ~io_inputBit | _GEN_5585; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5587 = i == 8'h2c ? _GEN_5586 : _GEN_5585; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5588 = io_inputBit ? 1'h0 : _GEN_5587; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5589 = i == 8'h2c ? _GEN_5588 : _GEN_5587; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5590 = io_inputBit | _GEN_5589; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5591 = i == 8'h51 ? _GEN_5590 : _GEN_5589; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5592 = ~io_inputBit ? 1'h0 : _GEN_5591; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5593 = i == 8'ha3 ? _GEN_5592 : _GEN_5591; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5594 = io_inputBit | _GEN_5593; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5596 = io_inputBit ? 1'h0 : _GEN_5171; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5597 = i == 8'h0 ? _GEN_5596 : _GEN_5171; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5598 = ~io_inputBit ? 1'h0 : _GEN_5597; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5599 = i == 8'h1 ? _GEN_5598 : _GEN_5597; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5600 = io_inputBit | _GEN_5599; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5601 = i == 8'h9 ? _GEN_5600 : _GEN_5599; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5602 = io_inputBit ? 1'h0 : _GEN_5601; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5603 = i == 8'h16 ? _GEN_5602 : _GEN_5601; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5604 = io_inputBit | _GEN_5603; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5605 = i == 8'h27 ? _GEN_5604 : _GEN_5603; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5606 = io_inputBit ? 1'h0 : _GEN_5605; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5607 = i == 8'h28 ? _GEN_5606 : _GEN_5605; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5608 = ~io_inputBit | _GEN_5607; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5609 = i == 8'h2b ? _GEN_5608 : _GEN_5607; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5610 = ~io_inputBit ? 1'h0 : _GEN_5609; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5611 = i == 8'h2c ? _GEN_5610 : _GEN_5609; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5612 = io_inputBit | _GEN_5611; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5613 = i == 8'h2c ? _GEN_5612 : _GEN_5611; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5614 = io_inputBit ? 1'h0 : _GEN_5613; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5615 = i == 8'h2d ? _GEN_5614 : _GEN_5613; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5616 = ~io_inputBit ? 1'h0 : _GEN_5615; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5617 = i == 8'h4f ? _GEN_5616 : _GEN_5615; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5618 = io_inputBit ? 1'h0 : _GEN_5617; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5619 = i == 8'h51 ? _GEN_5618 : _GEN_5617; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5620 = io_inputBit ? 1'h0 : _GEN_5619; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5621 = i == 8'h58 ? _GEN_5620 : _GEN_5619; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5622 = ~io_inputBit | _GEN_5621; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5623 = i == 8'h5b ? _GEN_5622 : _GEN_5621; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5624 = io_inputBit ? 1'h0 : _GEN_5623; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5625 = i == 8'h5b ? _GEN_5624 : _GEN_5623; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5626 = ~io_inputBit ? 1'h0 : _GEN_5625; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5627 = i == 8'ha0 ? _GEN_5626 : _GEN_5625; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5628 = io_inputBit | _GEN_5627; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5629 = i == 8'ha0 ? _GEN_5628 : _GEN_5627; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5630 = ~io_inputBit | _GEN_5629; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5631 = i == 8'ha3 ? _GEN_5630 : _GEN_5629; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5632 = io_inputBit ? 1'h0 : _GEN_5631; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5633 = i == 8'ha3 ? _GEN_5632 : _GEN_5631; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5634 = ~io_inputBit | _GEN_5633; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5635 = i == 8'hb1 ? _GEN_5634 : _GEN_5633; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5638 = io_inputBit ? 1'h0 : _GEN_5233; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5639 = i == 8'h0 ? _GEN_5638 : _GEN_5233; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5640 = ~io_inputBit ? 1'h0 : _GEN_5639; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5641 = i == 8'h1 ? _GEN_5640 : _GEN_5639; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5642 = io_inputBit ? 1'h0 : _GEN_5641; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5643 = i == 8'h9 ? _GEN_5642 : _GEN_5641; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5644 = io_inputBit ? 1'h0 : _GEN_5643; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5645 = i == 8'h16 ? _GEN_5644 : _GEN_5643; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5646 = io_inputBit | _GEN_5645; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5647 = i == 8'h28 ? _GEN_5646 : _GEN_5645; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5648 = ~io_inputBit ? 1'h0 : _GEN_5647; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5649 = i == 8'h2b ? _GEN_5648 : _GEN_5647; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5650 = ~io_inputBit | _GEN_5649; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5651 = i == 8'h4f ? _GEN_5650 : _GEN_5649; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5652 = ~io_inputBit ? 1'h0 : _GEN_5651; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5653 = i == 8'h50 ? _GEN_5652 : _GEN_5651; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5654 = io_inputBit | _GEN_5653; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5655 = i == 8'h50 ? _GEN_5654 : _GEN_5653; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5656 = io_inputBit ? 1'h0 : _GEN_5655; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5657 = i == 8'h51 ? _GEN_5656 : _GEN_5655; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5658 = io_inputBit | _GEN_5657; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5659 = i == 8'h58 ? _GEN_5658 : _GEN_5657; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5660 = io_inputBit ? 1'h0 : _GEN_5659; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5661 = i == 8'h59 ? _GEN_5660 : _GEN_5659; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5662 = ~io_inputBit | _GEN_5661; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5663 = i == 8'h5a ? _GEN_5662 : _GEN_5661; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5664 = ~io_inputBit ? 1'h0 : _GEN_5663; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5665 = i == 8'h5b ? _GEN_5664 : _GEN_5663; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5666 = io_inputBit | _GEN_5665; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5667 = i == 8'h5b ? _GEN_5666 : _GEN_5665; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5668 = io_inputBit ? 1'h0 : _GEN_5667; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5669 = i == 8'h5c ? _GEN_5668 : _GEN_5667; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5670 = ~io_inputBit | _GEN_5669; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5671 = i == 8'ha0 ? _GEN_5670 : _GEN_5669; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5672 = io_inputBit ? 1'h0 : _GEN_5671; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5673 = i == 8'ha0 ? _GEN_5672 : _GEN_5671; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5674 = ~io_inputBit | _GEN_5673; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5675 = i == 8'ha3 ? _GEN_5674 : _GEN_5673; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5676 = io_inputBit ? 1'h0 : _GEN_5675; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5677 = i == 8'ha3 ? _GEN_5676 : _GEN_5675; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5678 = ~io_inputBit ? 1'h0 : _GEN_5677; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5679 = i == 8'hb1 ? _GEN_5678 : _GEN_5677; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5680 = io_inputBit | _GEN_5679; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5681 = i == 8'hb1 ? _GEN_5680 : _GEN_5679; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5682 = ~io_inputBit | _GEN_5681; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5683 = i == 8'hb3 ? _GEN_5682 : _GEN_5681; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5684 = io_inputBit ? 1'h0 : _GEN_5683; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5685 = i == 8'hb3 ? _GEN_5684 : _GEN_5683; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5686 = ~io_inputBit | _GEN_5685; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5687 = i == 8'hb6 ? _GEN_5686 : _GEN_5685; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5688 = io_inputBit ? 1'h0 : _GEN_5687; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5689 = i == 8'hb6 ? _GEN_5688 : _GEN_5687; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5690 = ~io_inputBit | _GEN_5689; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5691 = i == 8'hb9 ? _GEN_5690 : _GEN_5689; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5694 = io_inputBit ? 1'h0 : _GEN_5313; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5695 = i == 8'h0 ? _GEN_5694 : _GEN_5313; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5696 = ~io_inputBit ? 1'h0 : _GEN_5695; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5697 = i == 8'h3 ? _GEN_5696 : _GEN_5695; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5698 = ~io_inputBit ? 1'h0 : _GEN_5697; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5699 = i == 8'h8 ? _GEN_5698 : _GEN_5697; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5700 = io_inputBit ? 1'h0 : _GEN_5699; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5701 = i == 8'h9 ? _GEN_5700 : _GEN_5699; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5702 = ~io_inputBit ? 1'h0 : _GEN_5701; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5703 = i == 8'h12 ? _GEN_5702 : _GEN_5701; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5704 = io_inputBit ? 1'h0 : _GEN_5703; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5705 = i == 8'h16 ? _GEN_5704 : _GEN_5703; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5706 = ~io_inputBit ? 1'h0 : _GEN_5705; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5707 = i == 8'h26 ? _GEN_5706 : _GEN_5705; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5708 = ~io_inputBit ? 1'h0 : _GEN_5707; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5709 = i == 8'h2b ? _GEN_5708 : _GEN_5707; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5710 = ~io_inputBit ? 1'h0 : _GEN_5709; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5711 = i == 8'h4e ? _GEN_5710 : _GEN_5709; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5712 = io_inputBit | _GEN_5711; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5713 = i == 8'h4e ? _GEN_5712 : _GEN_5711; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5714 = ~io_inputBit | _GEN_5713; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5715 = i == 8'h50 ? _GEN_5714 : _GEN_5713; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5716 = io_inputBit ? 1'h0 : _GEN_5715; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5717 = i == 8'h50 ? _GEN_5716 : _GEN_5715; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5718 = ~io_inputBit ? 1'h0 : _GEN_5717; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5719 = i == 8'h52 ? _GEN_5718 : _GEN_5717; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5720 = io_inputBit | _GEN_5719; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5721 = i == 8'h52 ? _GEN_5720 : _GEN_5719; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5722 = io_inputBit ? 1'h0 : _GEN_5721; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5723 = i == 8'h59 ? _GEN_5722 : _GEN_5721; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5724 = io_inputBit | _GEN_5723; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5725 = i == 8'h5b ? _GEN_5724 : _GEN_5723; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5726 = ~io_inputBit ? 1'h0 : _GEN_5725; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5727 = i == 8'h9f ? _GEN_5726 : _GEN_5725; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5728 = io_inputBit | _GEN_5727; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5729 = i == 8'h9f ? _GEN_5728 : _GEN_5727; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5730 = ~io_inputBit | _GEN_5729; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5731 = i == 8'ha0 ? _GEN_5730 : _GEN_5729; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5732 = io_inputBit ? 1'h0 : _GEN_5731; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5733 = i == 8'ha0 ? _GEN_5732 : _GEN_5731; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5734 = ~io_inputBit | _GEN_5733; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5735 = i == 8'ha3 ? _GEN_5734 : _GEN_5733; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5736 = io_inputBit ? 1'h0 : _GEN_5735; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5737 = i == 8'ha3 ? _GEN_5736 : _GEN_5735; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5738 = ~io_inputBit ? 1'h0 : _GEN_5737; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5739 = i == 8'ha4 ? _GEN_5738 : _GEN_5737; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5740 = io_inputBit | _GEN_5739; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5741 = i == 8'ha4 ? _GEN_5740 : _GEN_5739; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5742 = ~io_inputBit ? 1'h0 : _GEN_5741; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5743 = i == 8'hb1 ? _GEN_5742 : _GEN_5741; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5744 = io_inputBit | _GEN_5743; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5745 = i == 8'hb1 ? _GEN_5744 : _GEN_5743; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5746 = ~io_inputBit | _GEN_5745; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5747 = i == 8'hb2 ? _GEN_5746 : _GEN_5745; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5748 = io_inputBit ? 1'h0 : _GEN_5747; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5749 = i == 8'hb2 ? _GEN_5748 : _GEN_5747; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5750 = ~io_inputBit ? 1'h0 : _GEN_5749; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5751 = i == 8'hb3 ? _GEN_5750 : _GEN_5749; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5752 = io_inputBit | _GEN_5751; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5753 = i == 8'hb3 ? _GEN_5752 : _GEN_5751; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5754 = ~io_inputBit | _GEN_5753; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5755 = i == 8'hb5 ? _GEN_5754 : _GEN_5753; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5756 = io_inputBit ? 1'h0 : _GEN_5755; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5757 = i == 8'hb5 ? _GEN_5756 : _GEN_5755; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5758 = ~io_inputBit ? 1'h0 : _GEN_5757; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5759 = i == 8'hb6 ? _GEN_5758 : _GEN_5757; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5760 = io_inputBit | _GEN_5759; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5761 = i == 8'hb6 ? _GEN_5760 : _GEN_5759; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5762 = ~io_inputBit | _GEN_5761; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5763 = i == 8'hb7 ? _GEN_5762 : _GEN_5761; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5764 = io_inputBit ? 1'h0 : _GEN_5763; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5765 = i == 8'hb7 ? _GEN_5764 : _GEN_5763; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5766 = ~io_inputBit ? 1'h0 : _GEN_5765; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5767 = i == 8'hb9 ? _GEN_5766 : _GEN_5765; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5768 = io_inputBit | _GEN_5767; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5769 = i == 8'hb9 ? _GEN_5768 : _GEN_5767; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5770 = ~io_inputBit | _GEN_5769; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5771 = i == 8'hba ? _GEN_5770 : _GEN_5769; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5774 = io_inputBit ? 1'h0 : _GEN_5399; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5775 = i == 8'h0 ? _GEN_5774 : _GEN_5399; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5776 = ~io_inputBit ? 1'h0 : _GEN_5775; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5777 = i == 8'h3 ? _GEN_5776 : _GEN_5775; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5778 = ~io_inputBit ? 1'h0 : _GEN_5777; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5779 = i == 8'h8 ? _GEN_5778 : _GEN_5777; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5780 = io_inputBit | _GEN_5779; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5781 = i == 8'h9 ? _GEN_5780 : _GEN_5779; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5782 = ~io_inputBit ? 1'h0 : _GEN_5781; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5783 = i == 8'h12 ? _GEN_5782 : _GEN_5781; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5784 = io_inputBit ? 1'h0 : _GEN_5783; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5785 = i == 8'h16 ? _GEN_5784 : _GEN_5783; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5786 = ~io_inputBit ? 1'h0 : _GEN_5785; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5787 = i == 8'h26 ? _GEN_5786 : _GEN_5785; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5788 = ~io_inputBit | _GEN_5787; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5789 = i == 8'h2b ? _GEN_5788 : _GEN_5787; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5790 = ~io_inputBit | _GEN_5789; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5791 = i == 8'h58 ? _GEN_5790 : _GEN_5789; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5792 = ~io_inputBit ? 1'h0 : _GEN_5791; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5793 = i == 8'h59 ? _GEN_5792 : _GEN_5791; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5794 = ~io_inputBit | _GEN_5793; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5795 = i == 8'h5a ? _GEN_5794 : _GEN_5793; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5796 = ~io_inputBit ? 1'h0 : _GEN_5795; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5797 = i == 8'h5b ? _GEN_5796 : _GEN_5795; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5798 = ~io_inputBit | _GEN_5797; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5799 = i == 8'h5c ? _GEN_5798 : _GEN_5797; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5800 = ~io_inputBit ? 1'h0 : _GEN_5799; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5801 = i == 8'h9d ? _GEN_5800 : _GEN_5799; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5802 = io_inputBit | _GEN_5801; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5803 = i == 8'h9d ? _GEN_5802 : _GEN_5801; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5804 = ~io_inputBit ? 1'h0 : _GEN_5803; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5805 = i == 8'h9e ? _GEN_5804 : _GEN_5803; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5806 = io_inputBit | _GEN_5805; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5807 = i == 8'h9e ? _GEN_5806 : _GEN_5805; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5808 = ~io_inputBit | _GEN_5807; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5809 = i == 8'h9f ? _GEN_5808 : _GEN_5807; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5810 = io_inputBit ? 1'h0 : _GEN_5809; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5811 = i == 8'h9f ? _GEN_5810 : _GEN_5809; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5812 = ~io_inputBit | _GEN_5811; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5813 = i == 8'ha0 ? _GEN_5812 : _GEN_5811; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5814 = io_inputBit ? 1'h0 : _GEN_5813; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5815 = i == 8'ha0 ? _GEN_5814 : _GEN_5813; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5816 = ~io_inputBit ? 1'h0 : _GEN_5815; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5817 = i == 8'ha1 ? _GEN_5816 : _GEN_5815; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5818 = io_inputBit | _GEN_5817; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5819 = i == 8'ha1 ? _GEN_5818 : _GEN_5817; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5820 = ~io_inputBit ? 1'h0 : _GEN_5819; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5821 = i == 8'ha2 ? _GEN_5820 : _GEN_5819; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5822 = io_inputBit | _GEN_5821; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5823 = i == 8'ha2 ? _GEN_5822 : _GEN_5821; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5824 = ~io_inputBit | _GEN_5823; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5825 = i == 8'ha3 ? _GEN_5824 : _GEN_5823; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5826 = io_inputBit ? 1'h0 : _GEN_5825; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5827 = i == 8'ha3 ? _GEN_5826 : _GEN_5825; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5828 = ~io_inputBit | _GEN_5827; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5829 = i == 8'ha4 ? _GEN_5828 : _GEN_5827; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5830 = io_inputBit ? 1'h0 : _GEN_5829; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5831 = i == 8'ha4 ? _GEN_5830 : _GEN_5829; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5832 = ~io_inputBit ? 1'h0 : _GEN_5831; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5833 = i == 8'ha5 ? _GEN_5832 : _GEN_5831; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5834 = io_inputBit | _GEN_5833; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5835 = i == 8'ha5 ? _GEN_5834 : _GEN_5833; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5836 = ~io_inputBit ? 1'h0 : _GEN_5835; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5837 = i == 8'ha6 ? _GEN_5836 : _GEN_5835; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5838 = io_inputBit | _GEN_5837; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5839 = i == 8'ha6 ? _GEN_5838 : _GEN_5837; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5840 = ~io_inputBit ? 1'h0 : _GEN_5839; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5841 = i == 8'hb2 ? _GEN_5840 : _GEN_5839; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5842 = io_inputBit | _GEN_5841; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5843 = i == 8'hb2 ? _GEN_5842 : _GEN_5841; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5844 = ~io_inputBit | _GEN_5843; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5845 = i == 8'hb4 ? _GEN_5844 : _GEN_5843; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5846 = io_inputBit ? 1'h0 : _GEN_5845; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5847 = i == 8'hb4 ? _GEN_5846 : _GEN_5845; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5848 = ~io_inputBit ? 1'h0 : _GEN_5847; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5849 = i == 8'hb6 ? _GEN_5848 : _GEN_5847; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5850 = io_inputBit | _GEN_5849; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5851 = i == 8'hb6 ? _GEN_5850 : _GEN_5849; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5852 = ~io_inputBit | _GEN_5851; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5853 = i == 8'hb8 ? _GEN_5852 : _GEN_5851; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5854 = io_inputBit ? 1'h0 : _GEN_5853; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5855 = i == 8'hb8 ? _GEN_5854 : _GEN_5853; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5856 = ~io_inputBit ? 1'h0 : _GEN_5855; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5857 = i == 8'hba ? _GEN_5856 : _GEN_5855; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5858 = io_inputBit | _GEN_5857; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5860 = io_inputBit ? 1'h0 : _GEN_5475; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5861 = i == 8'h0 ? _GEN_5860 : _GEN_5475; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5862 = ~io_inputBit ? 1'h0 : _GEN_5861; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5863 = i == 8'h3 ? _GEN_5862 : _GEN_5861; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5864 = ~io_inputBit ? 1'h0 : _GEN_5863; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5865 = i == 8'h8 ? _GEN_5864 : _GEN_5863; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5866 = io_inputBit ? 1'h0 : _GEN_5865; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5867 = i == 8'h9 ? _GEN_5866 : _GEN_5865; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5868 = ~io_inputBit ? 1'h0 : _GEN_5867; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5869 = i == 8'h12 ? _GEN_5868 : _GEN_5867; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5870 = io_inputBit ? 1'h0 : _GEN_5869; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5871 = i == 8'h16 ? _GEN_5870 : _GEN_5869; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5872 = ~io_inputBit ? 1'h0 : _GEN_5871; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5873 = i == 8'h26 ? _GEN_5872 : _GEN_5871; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5874 = ~io_inputBit ? 1'h0 : _GEN_5873; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5875 = i == 8'h2b ? _GEN_5874 : _GEN_5873; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5876 = ~io_inputBit ? 1'h0 : _GEN_5875; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5877 = i == 8'h4e ? _GEN_5876 : _GEN_5875; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5878 = io_inputBit | _GEN_5877; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5879 = i == 8'h4e ? _GEN_5878 : _GEN_5877; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5880 = ~io_inputBit ? 1'h0 : _GEN_5879; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5881 = i == 8'h4f ? _GEN_5880 : _GEN_5879; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5882 = io_inputBit | _GEN_5881; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5883 = i == 8'h4f ? _GEN_5882 : _GEN_5881; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5884 = ~io_inputBit ? 1'h0 : _GEN_5883; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5885 = i == 8'h50 ? _GEN_5884 : _GEN_5883; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5886 = io_inputBit | _GEN_5885; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5887 = i == 8'h50 ? _GEN_5886 : _GEN_5885; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5888 = ~io_inputBit ? 1'h0 : _GEN_5887; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5889 = i == 8'h51 ? _GEN_5888 : _GEN_5887; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5890 = io_inputBit | _GEN_5889; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5891 = i == 8'h51 ? _GEN_5890 : _GEN_5889; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5892 = ~io_inputBit ? 1'h0 : _GEN_5891; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5893 = i == 8'h52 ? _GEN_5892 : _GEN_5891; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5894 = io_inputBit | _GEN_5893; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5895 = i == 8'h52 ? _GEN_5894 : _GEN_5893; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5896 = ~io_inputBit ? 1'h0 : _GEN_5895; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5897 = i == 8'hb1 ? _GEN_5896 : _GEN_5895; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5898 = io_inputBit | _GEN_5897; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5899 = i == 8'hb1 ? _GEN_5898 : _GEN_5897; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5900 = ~io_inputBit | _GEN_5899; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5901 = i == 8'hb2 ? _GEN_5900 : _GEN_5899; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5902 = io_inputBit ? 1'h0 : _GEN_5901; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5903 = i == 8'hb2 ? _GEN_5902 : _GEN_5901; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5904 = ~io_inputBit ? 1'h0 : _GEN_5903; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5905 = i == 8'hb3 ? _GEN_5904 : _GEN_5903; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5906 = io_inputBit | _GEN_5905; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5907 = i == 8'hb3 ? _GEN_5906 : _GEN_5905; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5908 = ~io_inputBit | _GEN_5907; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5909 = i == 8'hb4 ? _GEN_5908 : _GEN_5907; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5910 = io_inputBit ? 1'h0 : _GEN_5909; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5911 = i == 8'hb4 ? _GEN_5910 : _GEN_5909; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5912 = ~io_inputBit ? 1'h0 : _GEN_5911; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5913 = i == 8'hb5 ? _GEN_5912 : _GEN_5911; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5914 = io_inputBit | _GEN_5913; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5915 = i == 8'hb5 ? _GEN_5914 : _GEN_5913; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5916 = ~io_inputBit | _GEN_5915; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5917 = i == 8'hb6 ? _GEN_5916 : _GEN_5915; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5918 = io_inputBit ? 1'h0 : _GEN_5917; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5919 = i == 8'hb6 ? _GEN_5918 : _GEN_5917; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5920 = ~io_inputBit ? 1'h0 : _GEN_5919; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5921 = i == 8'hb7 ? _GEN_5920 : _GEN_5919; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5922 = io_inputBit | _GEN_5921; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5923 = i == 8'hb7 ? _GEN_5922 : _GEN_5921; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5924 = ~io_inputBit | _GEN_5923; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5925 = i == 8'hb8 ? _GEN_5924 : _GEN_5923; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5926 = io_inputBit ? 1'h0 : _GEN_5925; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5927 = i == 8'hb8 ? _GEN_5926 : _GEN_5925; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5928 = ~io_inputBit ? 1'h0 : _GEN_5927; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5929 = i == 8'hb9 ? _GEN_5928 : _GEN_5927; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5930 = io_inputBit | _GEN_5929; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5931 = i == 8'hb9 ? _GEN_5930 : _GEN_5929; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5932 = ~io_inputBit | _GEN_5931; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5933 = i == 8'hba ? _GEN_5932 : _GEN_5931; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5936 = io_inputBit ? 1'h0 : _GEN_5571; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5937 = i == 8'h0 ? _GEN_5936 : _GEN_5571; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5938 = ~io_inputBit ? 1'h0 : _GEN_5937; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5939 = i == 8'h3 ? _GEN_5938 : _GEN_5937; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5940 = ~io_inputBit ? 1'h0 : _GEN_5939; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5941 = i == 8'h8 ? _GEN_5940 : _GEN_5939; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5942 = io_inputBit ? 1'h0 : _GEN_5941; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5943 = i == 8'h9 ? _GEN_5942 : _GEN_5941; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5944 = ~io_inputBit ? 1'h0 : _GEN_5943; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5945 = i == 8'h12 ? _GEN_5944 : _GEN_5943; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5946 = io_inputBit ? 1'h0 : _GEN_5945; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5947 = i == 8'h16 ? _GEN_5946 : _GEN_5945; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5948 = ~io_inputBit ? 1'h0 : _GEN_5947; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5949 = i == 8'h26 ? _GEN_5948 : _GEN_5947; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5950 = ~io_inputBit ? 1'h0 : _GEN_5949; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5951 = i == 8'h2b ? _GEN_5950 : _GEN_5949; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5952 = ~io_inputBit ? 1'h0 : _GEN_5951; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5953 = i == 8'h9d ? _GEN_5952 : _GEN_5951; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5954 = io_inputBit | _GEN_5953; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5955 = i == 8'h9d ? _GEN_5954 : _GEN_5953; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5956 = ~io_inputBit ? 1'h0 : _GEN_5955; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5957 = i == 8'h9e ? _GEN_5956 : _GEN_5955; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5958 = io_inputBit | _GEN_5957; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5959 = i == 8'h9e ? _GEN_5958 : _GEN_5957; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5960 = ~io_inputBit ? 1'h0 : _GEN_5959; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5961 = i == 8'h9f ? _GEN_5960 : _GEN_5959; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5962 = io_inputBit | _GEN_5961; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5963 = i == 8'h9f ? _GEN_5962 : _GEN_5961; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5964 = ~io_inputBit ? 1'h0 : _GEN_5963; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5965 = i == 8'ha0 ? _GEN_5964 : _GEN_5963; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5966 = io_inputBit | _GEN_5965; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5967 = i == 8'ha0 ? _GEN_5966 : _GEN_5965; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5968 = ~io_inputBit ? 1'h0 : _GEN_5967; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5969 = i == 8'ha1 ? _GEN_5968 : _GEN_5967; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5970 = io_inputBit | _GEN_5969; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5971 = i == 8'ha1 ? _GEN_5970 : _GEN_5969; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5972 = ~io_inputBit ? 1'h0 : _GEN_5971; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5973 = i == 8'ha2 ? _GEN_5972 : _GEN_5971; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5974 = io_inputBit | _GEN_5973; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5975 = i == 8'ha2 ? _GEN_5974 : _GEN_5973; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5976 = ~io_inputBit ? 1'h0 : _GEN_5975; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5977 = i == 8'ha3 ? _GEN_5976 : _GEN_5975; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5978 = io_inputBit | _GEN_5977; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5979 = i == 8'ha3 ? _GEN_5978 : _GEN_5977; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5980 = ~io_inputBit ? 1'h0 : _GEN_5979; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5981 = i == 8'ha4 ? _GEN_5980 : _GEN_5979; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5982 = io_inputBit | _GEN_5981; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5983 = i == 8'ha4 ? _GEN_5982 : _GEN_5981; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5984 = ~io_inputBit ? 1'h0 : _GEN_5983; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5985 = i == 8'ha5 ? _GEN_5984 : _GEN_5983; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5986 = io_inputBit | _GEN_5985; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5987 = i == 8'ha5 ? _GEN_5986 : _GEN_5985; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5988 = ~io_inputBit ? 1'h0 : _GEN_5987; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5989 = i == 8'ha6 ? _GEN_5988 : _GEN_5987; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5990 = io_inputBit | _GEN_5989; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5991 = i == 8'ha6 ? _GEN_5990 : _GEN_5989; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5992 = ~io_inputBit ? 1'h0 : _GEN_5991; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5993 = i == 8'hb1 ? _GEN_5992 : _GEN_5991; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5994 = io_inputBit | _GEN_5993; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5995 = i == 8'hb1 ? _GEN_5994 : _GEN_5993; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5996 = ~io_inputBit ? 1'h0 : _GEN_5995; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5997 = i == 8'hb2 ? _GEN_5996 : _GEN_5995; // @[lut_mem_online.scala 235:34]
  wire  _GEN_5998 = io_inputBit | _GEN_5997; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_5999 = i == 8'hb2 ? _GEN_5998 : _GEN_5997; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6000 = ~io_inputBit ? 1'h0 : _GEN_5999; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6001 = i == 8'hb3 ? _GEN_6000 : _GEN_5999; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6002 = io_inputBit | _GEN_6001; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6003 = i == 8'hb3 ? _GEN_6002 : _GEN_6001; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6004 = ~io_inputBit ? 1'h0 : _GEN_6003; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6005 = i == 8'hb4 ? _GEN_6004 : _GEN_6003; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6006 = io_inputBit | _GEN_6005; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6007 = i == 8'hb4 ? _GEN_6006 : _GEN_6005; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6008 = ~io_inputBit ? 1'h0 : _GEN_6007; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6009 = i == 8'hb5 ? _GEN_6008 : _GEN_6007; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6010 = io_inputBit | _GEN_6009; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6011 = i == 8'hb5 ? _GEN_6010 : _GEN_6009; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6012 = ~io_inputBit ? 1'h0 : _GEN_6011; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6013 = i == 8'hb6 ? _GEN_6012 : _GEN_6011; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6014 = io_inputBit | _GEN_6013; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6015 = i == 8'hb6 ? _GEN_6014 : _GEN_6013; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6016 = ~io_inputBit ? 1'h0 : _GEN_6015; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6017 = i == 8'hb7 ? _GEN_6016 : _GEN_6015; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6018 = io_inputBit | _GEN_6017; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6019 = i == 8'hb7 ? _GEN_6018 : _GEN_6017; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6020 = ~io_inputBit ? 1'h0 : _GEN_6019; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6021 = i == 8'hb8 ? _GEN_6020 : _GEN_6019; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6022 = io_inputBit | _GEN_6021; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6023 = i == 8'hb8 ? _GEN_6022 : _GEN_6021; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6024 = ~io_inputBit ? 1'h0 : _GEN_6023; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6025 = i == 8'hb9 ? _GEN_6024 : _GEN_6023; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6026 = io_inputBit | _GEN_6025; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6027 = i == 8'hb9 ? _GEN_6026 : _GEN_6025; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6028 = ~io_inputBit ? 1'h0 : _GEN_6027; // @[lut_mem_online.scala 237:46 239:32]
  wire  _GEN_6029 = i == 8'hba ? _GEN_6028 : _GEN_6027; // @[lut_mem_online.scala 235:34]
  wire  _GEN_6030 = io_inputBit | _GEN_6029; // @[lut_mem_online.scala 237:46 239:32]
  wire  _T_6035 = counter < 5'h11; // @[lut_mem_online.scala 250:22]
  wire  _T_6036 = counter < 5'ha; // @[lut_mem_online.scala 255:24]
  wire  _T_6037 = counter >= 5'ha; // @[lut_mem_online.scala 258:30]
  wire [4:0] _outResult_T_1 = counter - 5'ha; // @[lut_mem_online.scala 260:41]
  wire  _GEN_6040 = 3'h1 == _outResult_T_1[2:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_6041 = 3'h2 == _outResult_T_1[2:0] ? buffer_2 : _GEN_6040; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_6042 = 3'h3 == _outResult_T_1[2:0] ? buffer_3 : _GEN_6041; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_6043 = 3'h4 == _outResult_T_1[2:0] ? buffer_4 : _GEN_6042; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_6044 = 3'h5 == _outResult_T_1[2:0] ? buffer_5 : _GEN_6043; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_6045 = 3'h6 == _outResult_T_1[2:0] ? buffer_6 : _GEN_6044; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_6046 = 3'h7 == _outResult_T_1[2:0] ? 1'h0 : _GEN_6045; // @[lut_mem_online.scala 260:{23,23}]
  wire  _T_6041 = ~reset; // @[lut_mem_online.scala 263:21]
  wire  _GEN_6048 = counter >= 5'ha ? _GEN_6046 : outResult; // @[lut_mem_online.scala 258:42 260:23 215:26]
  wire  _GEN_6050 = counter < 5'ha ? 1'h0 : _GEN_6048; // @[lut_mem_online.scala 255:35 257:23]
  wire  _T_6042 = i < 8'h7f; // @[lut_mem_online.scala 274:18]
  wire [9:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 284:24]
  wire [9:0] _i_T_2 = _i_T + 10'h1; // @[lut_mem_online.scala 284:28]
  wire [9:0] _i_T_5 = _i_T + 10'h2; // @[lut_mem_online.scala 286:28]
  wire [9:0] _GEN_6051 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 285:45 286:17 206:18]
  wire [9:0] _GEN_6052 = _T_10 ? _i_T_2 : _GEN_6051; // @[lut_mem_online.scala 283:39 284:17]
  wire  _T_6047 = i < 8'hff; // @[lut_mem_online.scala 289:24]
  wire [7:0] _GEN_6053 = i < 8'hff ? 8'hff : i; // @[lut_mem_online.scala 289:63 297:15 206:18]
  wire [9:0] _GEN_6054 = i < 8'h7f ? _GEN_6052 : {{2'd0}, _GEN_6053}; // @[lut_mem_online.scala 274:61]
  wire [4:0] _counter_T_1 = counter + 5'h1; // @[lut_mem_online.scala 300:30]
  wire  _GEN_6056 = counter < 5'h11 & _GEN_6050; // @[lut_mem_online.scala 250:52 304:21]
  wire [9:0] _GEN_6057 = counter < 5'h11 ? _GEN_6054 : {{2'd0}, i}; // @[lut_mem_online.scala 206:18 250:52]
  wire  _GEN_6080 = io_start & _GEN_6056; // @[lut_mem_online.scala 220:29 327:15]
  wire [9:0] _GEN_6081 = io_start ? _GEN_6057 : 10'h0; // @[lut_mem_online.scala 220:29 325:7]
  wire [9:0] _GEN_7910 = reset ? 10'h0 : _GEN_6081; // @[lut_mem_online.scala 206:{18,18}]
  wire  _GEN_7911 = io_start & _T_6035; // @[lut_mem_online.scala 263:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 334:16]
  always @(posedge clock) begin
    i <= _GEN_7910[7:0]; // @[lut_mem_online.scala 206:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'ha3) begin // @[lut_mem_online.scala 235:34]
          buffer_0 <= _GEN_5594;
        end else if (i == 8'ha3) begin // @[lut_mem_online.scala 235:34]
          buffer_0 <= _GEN_5592;
        end else begin
          buffer_0 <= _GEN_5591;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hb1) begin // @[lut_mem_online.scala 235:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 237:46]
            buffer_1 <= 1'h0; // @[lut_mem_online.scala 239:32]
          end else begin
            buffer_1 <= _GEN_5635;
          end
        end else begin
          buffer_1 <= _GEN_5635;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hb9) begin // @[lut_mem_online.scala 235:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 237:46]
            buffer_2 <= 1'h0; // @[lut_mem_online.scala 239:32]
          end else begin
            buffer_2 <= _GEN_5691;
          end
        end else begin
          buffer_2 <= _GEN_5691;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hba) begin // @[lut_mem_online.scala 235:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 237:46]
            buffer_3 <= 1'h0; // @[lut_mem_online.scala 239:32]
          end else begin
            buffer_3 <= _GEN_5771;
          end
        end else begin
          buffer_3 <= _GEN_5771;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hba) begin // @[lut_mem_online.scala 235:34]
          buffer_4 <= _GEN_5858;
        end else if (i == 8'hba) begin // @[lut_mem_online.scala 235:34]
          buffer_4 <= _GEN_5856;
        end else begin
          buffer_4 <= _GEN_5855;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hba) begin // @[lut_mem_online.scala 235:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 237:46]
            buffer_5 <= 1'h0; // @[lut_mem_online.scala 239:32]
          end else begin
            buffer_5 <= _GEN_5933;
          end
        end else begin
          buffer_5 <= _GEN_5933;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hba) begin // @[lut_mem_online.scala 235:34]
          buffer_6 <= _GEN_6030;
        end else if (i == 8'hba) begin // @[lut_mem_online.scala 235:34]
          buffer_6 <= _GEN_6028;
        end else begin
          buffer_6 <= _GEN_6027;
        end
      end
    end
    if (reset) begin // @[lut_mem_online.scala 212:24]
      counter <= 5'h0; // @[lut_mem_online.scala 212:24]
    end else if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h11) begin // @[lut_mem_online.scala 250:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 300:19]
      end
    end else begin
      counter <= 5'h0; // @[lut_mem_online.scala 326:13]
    end
    if (reset) begin // @[lut_mem_online.scala 215:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 215:26]
    end else begin
      outResult <= _GEN_6080;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_6035 & ~_T_6036 & _T_6037 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 263:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7911 & _T_6042 & _T_6041) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 277:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7911 & ~_T_6042 & _T_6047 & _T_6041) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 292:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
