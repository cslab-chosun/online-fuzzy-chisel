module RegularFuzzification(
  input        clock,
  input        reset,
  input        io_start,
  input  [9:0] io_inputs_0,
  input  [9:0] io_inputs_1,
  output       io_outResultValid,
  output [2:0] io_outResult
);
  wire [2:0] regMinVec_0_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_0_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_0_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_1_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_1_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_1_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_2_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_2_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_2_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_3_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_3_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_3_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_4_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_4_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_4_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_5_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_5_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_5_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_6_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_6_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_6_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_7_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_7_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_7_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_8_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_8_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_8_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_9_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_9_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_9_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_10_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_10_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_10_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_11_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_11_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_11_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_12_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_12_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_12_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_13_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_13_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_13_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_14_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_14_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_14_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_15_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_15_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_15_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_16_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_16_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_16_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_17_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_17_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_17_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_18_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_18_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_18_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_19_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_19_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_19_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_20_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_20_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_20_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_21_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_21_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_21_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_22_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_22_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_22_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_23_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_23_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_23_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_24_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [2:0] regMinVec_24_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_24_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire  regMaxVec_0_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_0_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_1_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_1_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_5; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_2_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_2_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_3_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_3_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_5; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_4_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_4_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  outResult_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  outResult_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  reg [2:0] regLutResultsVec_0; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_1; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_2; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_3; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_4; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_5; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_6; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_7; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_8; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_9; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regMinVec_0; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_1; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_2; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_3; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_4; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_5; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_6; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_7; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_8; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_9; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_10; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_11; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_12; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_13; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_14; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_15; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_16; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_17; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_18; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_19; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_20; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_21; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_22; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_23; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_24; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMaxVec_0; // @[regular_fuzzification.scala 159:22]
  reg [2:0] regMaxVec_1; // @[regular_fuzzification.scala 159:22]
  reg [2:0] regMaxVec_2; // @[regular_fuzzification.scala 159:22]
  reg [2:0] regMaxVec_3; // @[regular_fuzzification.scala 159:22]
  reg [2:0] regMaxVec_4; // @[regular_fuzzification.scala 159:22]
  wire [6:0] _GEN_21 = 8'h15 == io_inputs_0[7:0] ? 7'h5f : 7'h64; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_22 = 8'h16 == io_inputs_0[7:0] ? 7'h5a : _GEN_21; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_23 = 8'h17 == io_inputs_0[7:0] ? 7'h55 : _GEN_22; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_24 = 8'h18 == io_inputs_0[7:0] ? 7'h50 : _GEN_23; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_25 = 8'h19 == io_inputs_0[7:0] ? 7'h4b : _GEN_24; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_26 = 8'h1a == io_inputs_0[7:0] ? 7'h46 : _GEN_25; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_27 = 8'h1b == io_inputs_0[7:0] ? 7'h41 : _GEN_26; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_28 = 8'h1c == io_inputs_0[7:0] ? 7'h3c : _GEN_27; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_29 = 8'h1d == io_inputs_0[7:0] ? 7'h37 : _GEN_28; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_30 = 8'h1e == io_inputs_0[7:0] ? 7'h32 : _GEN_29; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_31 = 8'h1f == io_inputs_0[7:0] ? 7'h2d : _GEN_30; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_32 = 8'h20 == io_inputs_0[7:0] ? 7'h28 : _GEN_31; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_33 = 8'h21 == io_inputs_0[7:0] ? 7'h23 : _GEN_32; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_34 = 8'h22 == io_inputs_0[7:0] ? 7'h1e : _GEN_33; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_35 = 8'h23 == io_inputs_0[7:0] ? 7'h19 : _GEN_34; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_36 = 8'h24 == io_inputs_0[7:0] ? 7'h14 : _GEN_35; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_37 = 8'h25 == io_inputs_0[7:0] ? 7'hf : _GEN_36; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_38 = 8'h26 == io_inputs_0[7:0] ? 7'ha : _GEN_37; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_39 = 8'h27 == io_inputs_0[7:0] ? 7'h5 : _GEN_38; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_40 = 8'h28 == io_inputs_0[7:0] ? 7'h0 : _GEN_39; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_41 = 8'h29 == io_inputs_0[7:0] ? 7'h0 : _GEN_40; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_42 = 8'h2a == io_inputs_0[7:0] ? 7'h0 : _GEN_41; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_43 = 8'h2b == io_inputs_0[7:0] ? 7'h0 : _GEN_42; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_44 = 8'h2c == io_inputs_0[7:0] ? 7'h0 : _GEN_43; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_45 = 8'h2d == io_inputs_0[7:0] ? 7'h0 : _GEN_44; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_46 = 8'h2e == io_inputs_0[7:0] ? 7'h0 : _GEN_45; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_47 = 8'h2f == io_inputs_0[7:0] ? 7'h0 : _GEN_46; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_48 = 8'h30 == io_inputs_0[7:0] ? 7'h0 : _GEN_47; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_49 = 8'h31 == io_inputs_0[7:0] ? 7'h0 : _GEN_48; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_50 = 8'h32 == io_inputs_0[7:0] ? 7'h0 : _GEN_49; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_51 = 8'h33 == io_inputs_0[7:0] ? 7'h0 : _GEN_50; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_52 = 8'h34 == io_inputs_0[7:0] ? 7'h0 : _GEN_51; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_53 = 8'h35 == io_inputs_0[7:0] ? 7'h0 : _GEN_52; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_54 = 8'h36 == io_inputs_0[7:0] ? 7'h0 : _GEN_53; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_55 = 8'h37 == io_inputs_0[7:0] ? 7'h0 : _GEN_54; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_56 = 8'h38 == io_inputs_0[7:0] ? 7'h0 : _GEN_55; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_57 = 8'h39 == io_inputs_0[7:0] ? 7'h0 : _GEN_56; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_58 = 8'h3a == io_inputs_0[7:0] ? 7'h0 : _GEN_57; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_59 = 8'h3b == io_inputs_0[7:0] ? 7'h0 : _GEN_58; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_60 = 8'h3c == io_inputs_0[7:0] ? 7'h0 : _GEN_59; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_61 = 8'h3d == io_inputs_0[7:0] ? 7'h0 : _GEN_60; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_62 = 8'h3e == io_inputs_0[7:0] ? 7'h0 : _GEN_61; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_63 = 8'h3f == io_inputs_0[7:0] ? 7'h0 : _GEN_62; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_64 = 8'h40 == io_inputs_0[7:0] ? 7'h0 : _GEN_63; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_65 = 8'h41 == io_inputs_0[7:0] ? 7'h0 : _GEN_64; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_66 = 8'h42 == io_inputs_0[7:0] ? 7'h0 : _GEN_65; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_67 = 8'h43 == io_inputs_0[7:0] ? 7'h0 : _GEN_66; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_68 = 8'h44 == io_inputs_0[7:0] ? 7'h0 : _GEN_67; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_69 = 8'h45 == io_inputs_0[7:0] ? 7'h0 : _GEN_68; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_70 = 8'h46 == io_inputs_0[7:0] ? 7'h0 : _GEN_69; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_71 = 8'h47 == io_inputs_0[7:0] ? 7'h0 : _GEN_70; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_72 = 8'h48 == io_inputs_0[7:0] ? 7'h0 : _GEN_71; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_73 = 8'h49 == io_inputs_0[7:0] ? 7'h0 : _GEN_72; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_74 = 8'h4a == io_inputs_0[7:0] ? 7'h0 : _GEN_73; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_75 = 8'h4b == io_inputs_0[7:0] ? 7'h0 : _GEN_74; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_76 = 8'h4c == io_inputs_0[7:0] ? 7'h0 : _GEN_75; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_77 = 8'h4d == io_inputs_0[7:0] ? 7'h0 : _GEN_76; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_78 = 8'h4e == io_inputs_0[7:0] ? 7'h0 : _GEN_77; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_79 = 8'h4f == io_inputs_0[7:0] ? 7'h0 : _GEN_78; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_80 = 8'h50 == io_inputs_0[7:0] ? 7'h0 : _GEN_79; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_81 = 8'h51 == io_inputs_0[7:0] ? 7'h0 : _GEN_80; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_82 = 8'h52 == io_inputs_0[7:0] ? 7'h0 : _GEN_81; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_83 = 8'h53 == io_inputs_0[7:0] ? 7'h0 : _GEN_82; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_84 = 8'h54 == io_inputs_0[7:0] ? 7'h0 : _GEN_83; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_85 = 8'h55 == io_inputs_0[7:0] ? 7'h0 : _GEN_84; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_86 = 8'h56 == io_inputs_0[7:0] ? 7'h0 : _GEN_85; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_87 = 8'h57 == io_inputs_0[7:0] ? 7'h0 : _GEN_86; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_88 = 8'h58 == io_inputs_0[7:0] ? 7'h0 : _GEN_87; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_89 = 8'h59 == io_inputs_0[7:0] ? 7'h0 : _GEN_88; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_90 = 8'h5a == io_inputs_0[7:0] ? 7'h0 : _GEN_89; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_91 = 8'h5b == io_inputs_0[7:0] ? 7'h0 : _GEN_90; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_92 = 8'h5c == io_inputs_0[7:0] ? 7'h0 : _GEN_91; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_93 = 8'h5d == io_inputs_0[7:0] ? 7'h0 : _GEN_92; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_94 = 8'h5e == io_inputs_0[7:0] ? 7'h0 : _GEN_93; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_95 = 8'h5f == io_inputs_0[7:0] ? 7'h0 : _GEN_94; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_96 = 8'h60 == io_inputs_0[7:0] ? 7'h0 : _GEN_95; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_97 = 8'h61 == io_inputs_0[7:0] ? 7'h0 : _GEN_96; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_98 = 8'h62 == io_inputs_0[7:0] ? 7'h0 : _GEN_97; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_99 = 8'h63 == io_inputs_0[7:0] ? 7'h0 : _GEN_98; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_100 = 8'h64 == io_inputs_0[7:0] ? 7'h0 : _GEN_99; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_101 = 8'h65 == io_inputs_0[7:0] ? 7'h0 : _GEN_100; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_102 = 8'h66 == io_inputs_0[7:0] ? 7'h0 : _GEN_101; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_103 = 8'h67 == io_inputs_0[7:0] ? 7'h0 : _GEN_102; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_104 = 8'h68 == io_inputs_0[7:0] ? 7'h0 : _GEN_103; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_105 = 8'h69 == io_inputs_0[7:0] ? 7'h0 : _GEN_104; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_106 = 8'h6a == io_inputs_0[7:0] ? 7'h0 : _GEN_105; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_107 = 8'h6b == io_inputs_0[7:0] ? 7'h0 : _GEN_106; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_108 = 8'h6c == io_inputs_0[7:0] ? 7'h0 : _GEN_107; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_109 = 8'h6d == io_inputs_0[7:0] ? 7'h0 : _GEN_108; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_110 = 8'h6e == io_inputs_0[7:0] ? 7'h0 : _GEN_109; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_111 = 8'h6f == io_inputs_0[7:0] ? 7'h0 : _GEN_110; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_112 = 8'h70 == io_inputs_0[7:0] ? 7'h0 : _GEN_111; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_113 = 8'h71 == io_inputs_0[7:0] ? 7'h0 : _GEN_112; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_114 = 8'h72 == io_inputs_0[7:0] ? 7'h0 : _GEN_113; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_115 = 8'h73 == io_inputs_0[7:0] ? 7'h0 : _GEN_114; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_116 = 8'h74 == io_inputs_0[7:0] ? 7'h0 : _GEN_115; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_117 = 8'h75 == io_inputs_0[7:0] ? 7'h0 : _GEN_116; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_118 = 8'h76 == io_inputs_0[7:0] ? 7'h0 : _GEN_117; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_119 = 8'h77 == io_inputs_0[7:0] ? 7'h0 : _GEN_118; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_120 = 8'h78 == io_inputs_0[7:0] ? 7'h0 : _GEN_119; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_121 = 8'h79 == io_inputs_0[7:0] ? 7'h0 : _GEN_120; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_122 = 8'h7a == io_inputs_0[7:0] ? 7'h0 : _GEN_121; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_123 = 8'h7b == io_inputs_0[7:0] ? 7'h0 : _GEN_122; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_124 = 8'h7c == io_inputs_0[7:0] ? 7'h0 : _GEN_123; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_125 = 8'h7d == io_inputs_0[7:0] ? 7'h0 : _GEN_124; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_126 = 8'h7e == io_inputs_0[7:0] ? 7'h0 : _GEN_125; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_127 = 8'h7f == io_inputs_0[7:0] ? 7'h0 : _GEN_126; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_128 = 8'h80 == io_inputs_0[7:0] ? 7'h0 : _GEN_127; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_129 = 8'h81 == io_inputs_0[7:0] ? 7'h0 : _GEN_128; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_130 = 8'h82 == io_inputs_0[7:0] ? 7'h0 : _GEN_129; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_131 = 8'h83 == io_inputs_0[7:0] ? 7'h0 : _GEN_130; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_132 = 8'h84 == io_inputs_0[7:0] ? 7'h0 : _GEN_131; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_133 = 8'h85 == io_inputs_0[7:0] ? 7'h0 : _GEN_132; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_134 = 8'h86 == io_inputs_0[7:0] ? 7'h0 : _GEN_133; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_135 = 8'h87 == io_inputs_0[7:0] ? 7'h0 : _GEN_134; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_136 = 8'h88 == io_inputs_0[7:0] ? 7'h0 : _GEN_135; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_137 = 8'h89 == io_inputs_0[7:0] ? 7'h0 : _GEN_136; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_138 = 8'h8a == io_inputs_0[7:0] ? 7'h0 : _GEN_137; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_139 = 8'h8b == io_inputs_0[7:0] ? 7'h0 : _GEN_138; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_140 = 8'h8c == io_inputs_0[7:0] ? 7'h0 : _GEN_139; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_141 = 8'h8d == io_inputs_0[7:0] ? 7'h0 : _GEN_140; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_142 = 8'h8e == io_inputs_0[7:0] ? 7'h0 : _GEN_141; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_143 = 8'h8f == io_inputs_0[7:0] ? 7'h0 : _GEN_142; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_144 = 8'h90 == io_inputs_0[7:0] ? 7'h0 : _GEN_143; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_145 = 8'h91 == io_inputs_0[7:0] ? 7'h0 : _GEN_144; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_146 = 8'h92 == io_inputs_0[7:0] ? 7'h0 : _GEN_145; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_147 = 8'h93 == io_inputs_0[7:0] ? 7'h0 : _GEN_146; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_148 = 8'h94 == io_inputs_0[7:0] ? 7'h0 : _GEN_147; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_149 = 8'h95 == io_inputs_0[7:0] ? 7'h0 : _GEN_148; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_150 = 8'h96 == io_inputs_0[7:0] ? 7'h0 : _GEN_149; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_151 = 8'h97 == io_inputs_0[7:0] ? 7'h0 : _GEN_150; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_152 = 8'h98 == io_inputs_0[7:0] ? 7'h0 : _GEN_151; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_153 = 8'h99 == io_inputs_0[7:0] ? 7'h0 : _GEN_152; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_154 = 8'h9a == io_inputs_0[7:0] ? 7'h0 : _GEN_153; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_155 = 8'h9b == io_inputs_0[7:0] ? 7'h0 : _GEN_154; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_156 = 8'h9c == io_inputs_0[7:0] ? 7'h0 : _GEN_155; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_157 = 8'h9d == io_inputs_0[7:0] ? 7'h0 : _GEN_156; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_158 = 8'h9e == io_inputs_0[7:0] ? 7'h0 : _GEN_157; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_159 = 8'h9f == io_inputs_0[7:0] ? 7'h0 : _GEN_158; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_160 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_159; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_161 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_160; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_162 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_161; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_163 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_162; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_164 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_163; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_165 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_164; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_166 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_167 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_168 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_169 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_170 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_171 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_172 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_173 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_174 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_175 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_176 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_177 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_178 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_179 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_180 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_181 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_182 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_183 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_184 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_185 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_186 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_187 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_188 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_189 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_190 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_191 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_192 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_193 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_194 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_195 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_196 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_197 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_198 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_199 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_200 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_201 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_202 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_203 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_204 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_205 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_206 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_207 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_208 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_209 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_210 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_211 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_212 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_213 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_214 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_215 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_216 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_217 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_218 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_219 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_220 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_221 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_222 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_223 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_224 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_225 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_226 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_227 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_228 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_229 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_230 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_231 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_232 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_233 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_234 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_235 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_236 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_237 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_238 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_239 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_240 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_241 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_242 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_243 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_244 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_245 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_246 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_247 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_248 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_249 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_250 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_251 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_252 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_253 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_254 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_255 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_277 = 8'h15 == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_278 = 8'h16 == io_inputs_0[7:0] ? 7'ha : _GEN_277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_279 = 8'h17 == io_inputs_0[7:0] ? 7'hf : _GEN_278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_280 = 8'h18 == io_inputs_0[7:0] ? 7'h14 : _GEN_279; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_281 = 8'h19 == io_inputs_0[7:0] ? 7'h19 : _GEN_280; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_282 = 8'h1a == io_inputs_0[7:0] ? 7'h1e : _GEN_281; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_283 = 8'h1b == io_inputs_0[7:0] ? 7'h23 : _GEN_282; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_284 = 8'h1c == io_inputs_0[7:0] ? 7'h28 : _GEN_283; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_285 = 8'h1d == io_inputs_0[7:0] ? 7'h2d : _GEN_284; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_286 = 8'h1e == io_inputs_0[7:0] ? 7'h32 : _GEN_285; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_287 = 8'h1f == io_inputs_0[7:0] ? 7'h37 : _GEN_286; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_288 = 8'h20 == io_inputs_0[7:0] ? 7'h3c : _GEN_287; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_289 = 8'h21 == io_inputs_0[7:0] ? 7'h41 : _GEN_288; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_290 = 8'h22 == io_inputs_0[7:0] ? 7'h46 : _GEN_289; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_291 = 8'h23 == io_inputs_0[7:0] ? 7'h4b : _GEN_290; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_292 = 8'h24 == io_inputs_0[7:0] ? 7'h50 : _GEN_291; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_293 = 8'h25 == io_inputs_0[7:0] ? 7'h55 : _GEN_292; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_294 = 8'h26 == io_inputs_0[7:0] ? 7'h5a : _GEN_293; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_295 = 8'h27 == io_inputs_0[7:0] ? 7'h5f : _GEN_294; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_296 = 8'h28 == io_inputs_0[7:0] ? 7'h64 : _GEN_295; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_297 = 8'h29 == io_inputs_0[7:0] ? 7'h64 : _GEN_296; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_298 = 8'h2a == io_inputs_0[7:0] ? 7'h64 : _GEN_297; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_299 = 8'h2b == io_inputs_0[7:0] ? 7'h64 : _GEN_298; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_300 = 8'h2c == io_inputs_0[7:0] ? 7'h64 : _GEN_299; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_301 = 8'h2d == io_inputs_0[7:0] ? 7'h64 : _GEN_300; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_302 = 8'h2e == io_inputs_0[7:0] ? 7'h64 : _GEN_301; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_303 = 8'h2f == io_inputs_0[7:0] ? 7'h64 : _GEN_302; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_304 = 8'h30 == io_inputs_0[7:0] ? 7'h64 : _GEN_303; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_305 = 8'h31 == io_inputs_0[7:0] ? 7'h64 : _GEN_304; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_306 = 8'h32 == io_inputs_0[7:0] ? 7'h64 : _GEN_305; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_307 = 8'h33 == io_inputs_0[7:0] ? 7'h64 : _GEN_306; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_308 = 8'h34 == io_inputs_0[7:0] ? 7'h64 : _GEN_307; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_309 = 8'h35 == io_inputs_0[7:0] ? 7'h64 : _GEN_308; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_310 = 8'h36 == io_inputs_0[7:0] ? 7'h64 : _GEN_309; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_311 = 8'h37 == io_inputs_0[7:0] ? 7'h64 : _GEN_310; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_312 = 8'h38 == io_inputs_0[7:0] ? 7'h64 : _GEN_311; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_313 = 8'h39 == io_inputs_0[7:0] ? 7'h64 : _GEN_312; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_314 = 8'h3a == io_inputs_0[7:0] ? 7'h64 : _GEN_313; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_315 = 8'h3b == io_inputs_0[7:0] ? 7'h64 : _GEN_314; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_316 = 8'h3c == io_inputs_0[7:0] ? 7'h64 : _GEN_315; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_317 = 8'h3d == io_inputs_0[7:0] ? 7'h5f : _GEN_316; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_318 = 8'h3e == io_inputs_0[7:0] ? 7'h5a : _GEN_317; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_319 = 8'h3f == io_inputs_0[7:0] ? 7'h55 : _GEN_318; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_320 = 8'h40 == io_inputs_0[7:0] ? 7'h50 : _GEN_319; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_321 = 8'h41 == io_inputs_0[7:0] ? 7'h4b : _GEN_320; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_322 = 8'h42 == io_inputs_0[7:0] ? 7'h46 : _GEN_321; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_323 = 8'h43 == io_inputs_0[7:0] ? 7'h41 : _GEN_322; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_324 = 8'h44 == io_inputs_0[7:0] ? 7'h3c : _GEN_323; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_325 = 8'h45 == io_inputs_0[7:0] ? 7'h37 : _GEN_324; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_326 = 8'h46 == io_inputs_0[7:0] ? 7'h32 : _GEN_325; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_327 = 8'h47 == io_inputs_0[7:0] ? 7'h2d : _GEN_326; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_328 = 8'h48 == io_inputs_0[7:0] ? 7'h28 : _GEN_327; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_329 = 8'h49 == io_inputs_0[7:0] ? 7'h23 : _GEN_328; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_330 = 8'h4a == io_inputs_0[7:0] ? 7'h1e : _GEN_329; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_331 = 8'h4b == io_inputs_0[7:0] ? 7'h19 : _GEN_330; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_332 = 8'h4c == io_inputs_0[7:0] ? 7'h14 : _GEN_331; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_333 = 8'h4d == io_inputs_0[7:0] ? 7'hf : _GEN_332; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_334 = 8'h4e == io_inputs_0[7:0] ? 7'ha : _GEN_333; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_335 = 8'h4f == io_inputs_0[7:0] ? 7'h5 : _GEN_334; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_336 = 8'h50 == io_inputs_0[7:0] ? 7'h0 : _GEN_335; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_337 = 8'h51 == io_inputs_0[7:0] ? 7'h0 : _GEN_336; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_338 = 8'h52 == io_inputs_0[7:0] ? 7'h0 : _GEN_337; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_339 = 8'h53 == io_inputs_0[7:0] ? 7'h0 : _GEN_338; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_340 = 8'h54 == io_inputs_0[7:0] ? 7'h0 : _GEN_339; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_341 = 8'h55 == io_inputs_0[7:0] ? 7'h0 : _GEN_340; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_342 = 8'h56 == io_inputs_0[7:0] ? 7'h0 : _GEN_341; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_343 = 8'h57 == io_inputs_0[7:0] ? 7'h0 : _GEN_342; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_344 = 8'h58 == io_inputs_0[7:0] ? 7'h0 : _GEN_343; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_345 = 8'h59 == io_inputs_0[7:0] ? 7'h0 : _GEN_344; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_346 = 8'h5a == io_inputs_0[7:0] ? 7'h0 : _GEN_345; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_347 = 8'h5b == io_inputs_0[7:0] ? 7'h0 : _GEN_346; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_348 = 8'h5c == io_inputs_0[7:0] ? 7'h0 : _GEN_347; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_349 = 8'h5d == io_inputs_0[7:0] ? 7'h0 : _GEN_348; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_350 = 8'h5e == io_inputs_0[7:0] ? 7'h0 : _GEN_349; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_351 = 8'h5f == io_inputs_0[7:0] ? 7'h0 : _GEN_350; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_352 = 8'h60 == io_inputs_0[7:0] ? 7'h0 : _GEN_351; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_353 = 8'h61 == io_inputs_0[7:0] ? 7'h0 : _GEN_352; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_354 = 8'h62 == io_inputs_0[7:0] ? 7'h0 : _GEN_353; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_355 = 8'h63 == io_inputs_0[7:0] ? 7'h0 : _GEN_354; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_356 = 8'h64 == io_inputs_0[7:0] ? 7'h0 : _GEN_355; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_357 = 8'h65 == io_inputs_0[7:0] ? 7'h0 : _GEN_356; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_358 = 8'h66 == io_inputs_0[7:0] ? 7'h0 : _GEN_357; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_359 = 8'h67 == io_inputs_0[7:0] ? 7'h0 : _GEN_358; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_360 = 8'h68 == io_inputs_0[7:0] ? 7'h0 : _GEN_359; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_361 = 8'h69 == io_inputs_0[7:0] ? 7'h0 : _GEN_360; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_362 = 8'h6a == io_inputs_0[7:0] ? 7'h0 : _GEN_361; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_363 = 8'h6b == io_inputs_0[7:0] ? 7'h0 : _GEN_362; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_364 = 8'h6c == io_inputs_0[7:0] ? 7'h0 : _GEN_363; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_365 = 8'h6d == io_inputs_0[7:0] ? 7'h0 : _GEN_364; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_366 = 8'h6e == io_inputs_0[7:0] ? 7'h0 : _GEN_365; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_367 = 8'h6f == io_inputs_0[7:0] ? 7'h0 : _GEN_366; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_368 = 8'h70 == io_inputs_0[7:0] ? 7'h0 : _GEN_367; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_369 = 8'h71 == io_inputs_0[7:0] ? 7'h0 : _GEN_368; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_370 = 8'h72 == io_inputs_0[7:0] ? 7'h0 : _GEN_369; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_371 = 8'h73 == io_inputs_0[7:0] ? 7'h0 : _GEN_370; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_372 = 8'h74 == io_inputs_0[7:0] ? 7'h0 : _GEN_371; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_373 = 8'h75 == io_inputs_0[7:0] ? 7'h0 : _GEN_372; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_374 = 8'h76 == io_inputs_0[7:0] ? 7'h0 : _GEN_373; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_375 = 8'h77 == io_inputs_0[7:0] ? 7'h0 : _GEN_374; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_376 = 8'h78 == io_inputs_0[7:0] ? 7'h0 : _GEN_375; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_377 = 8'h79 == io_inputs_0[7:0] ? 7'h0 : _GEN_376; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_378 = 8'h7a == io_inputs_0[7:0] ? 7'h0 : _GEN_377; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_379 = 8'h7b == io_inputs_0[7:0] ? 7'h0 : _GEN_378; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_380 = 8'h7c == io_inputs_0[7:0] ? 7'h0 : _GEN_379; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_381 = 8'h7d == io_inputs_0[7:0] ? 7'h0 : _GEN_380; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_382 = 8'h7e == io_inputs_0[7:0] ? 7'h0 : _GEN_381; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_383 = 8'h7f == io_inputs_0[7:0] ? 7'h0 : _GEN_382; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_384 = 8'h80 == io_inputs_0[7:0] ? 7'h0 : _GEN_383; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_385 = 8'h81 == io_inputs_0[7:0] ? 7'h0 : _GEN_384; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_386 = 8'h82 == io_inputs_0[7:0] ? 7'h0 : _GEN_385; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_387 = 8'h83 == io_inputs_0[7:0] ? 7'h0 : _GEN_386; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_388 = 8'h84 == io_inputs_0[7:0] ? 7'h0 : _GEN_387; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_389 = 8'h85 == io_inputs_0[7:0] ? 7'h0 : _GEN_388; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_390 = 8'h86 == io_inputs_0[7:0] ? 7'h0 : _GEN_389; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_391 = 8'h87 == io_inputs_0[7:0] ? 7'h0 : _GEN_390; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_392 = 8'h88 == io_inputs_0[7:0] ? 7'h0 : _GEN_391; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_393 = 8'h89 == io_inputs_0[7:0] ? 7'h0 : _GEN_392; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_394 = 8'h8a == io_inputs_0[7:0] ? 7'h0 : _GEN_393; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_395 = 8'h8b == io_inputs_0[7:0] ? 7'h0 : _GEN_394; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_396 = 8'h8c == io_inputs_0[7:0] ? 7'h0 : _GEN_395; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_397 = 8'h8d == io_inputs_0[7:0] ? 7'h0 : _GEN_396; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_398 = 8'h8e == io_inputs_0[7:0] ? 7'h0 : _GEN_397; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_399 = 8'h8f == io_inputs_0[7:0] ? 7'h0 : _GEN_398; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_400 = 8'h90 == io_inputs_0[7:0] ? 7'h0 : _GEN_399; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_401 = 8'h91 == io_inputs_0[7:0] ? 7'h0 : _GEN_400; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_402 = 8'h92 == io_inputs_0[7:0] ? 7'h0 : _GEN_401; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_403 = 8'h93 == io_inputs_0[7:0] ? 7'h0 : _GEN_402; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_404 = 8'h94 == io_inputs_0[7:0] ? 7'h0 : _GEN_403; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_405 = 8'h95 == io_inputs_0[7:0] ? 7'h0 : _GEN_404; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_406 = 8'h96 == io_inputs_0[7:0] ? 7'h0 : _GEN_405; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_407 = 8'h97 == io_inputs_0[7:0] ? 7'h0 : _GEN_406; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_408 = 8'h98 == io_inputs_0[7:0] ? 7'h0 : _GEN_407; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_409 = 8'h99 == io_inputs_0[7:0] ? 7'h0 : _GEN_408; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_410 = 8'h9a == io_inputs_0[7:0] ? 7'h0 : _GEN_409; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_411 = 8'h9b == io_inputs_0[7:0] ? 7'h0 : _GEN_410; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_412 = 8'h9c == io_inputs_0[7:0] ? 7'h0 : _GEN_411; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_413 = 8'h9d == io_inputs_0[7:0] ? 7'h0 : _GEN_412; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_414 = 8'h9e == io_inputs_0[7:0] ? 7'h0 : _GEN_413; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_415 = 8'h9f == io_inputs_0[7:0] ? 7'h0 : _GEN_414; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_416 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_415; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_417 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_416; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_418 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_417; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_419 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_418; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_420 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_419; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_421 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_420; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_422 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_421; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_423 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_422; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_424 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_423; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_425 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_424; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_426 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_425; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_427 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_426; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_428 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_427; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_429 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_428; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_430 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_429; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_431 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_430; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_432 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_431; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_433 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_432; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_434 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_433; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_435 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_434; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_436 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_435; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_437 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_436; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_438 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_437; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_439 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_438; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_440 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_439; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_441 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_440; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_442 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_441; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_443 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_442; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_444 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_443; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_445 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_444; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_446 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_445; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_447 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_446; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_448 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_447; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_449 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_448; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_450 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_449; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_451 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_450; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_452 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_451; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_453 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_452; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_454 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_453; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_455 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_454; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_456 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_455; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_457 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_456; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_458 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_457; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_459 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_458; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_460 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_459; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_461 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_460; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_462 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_461; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_463 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_462; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_464 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_463; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_465 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_464; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_466 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_465; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_467 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_466; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_468 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_467; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_469 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_468; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_470 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_469; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_471 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_470; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_472 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_471; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_473 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_472; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_474 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_473; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_475 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_474; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_476 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_475; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_477 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_476; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_478 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_477; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_479 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_478; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_480 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_479; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_481 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_480; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_482 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_481; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_483 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_482; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_484 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_483; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_485 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_484; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_486 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_485; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_487 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_486; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_488 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_487; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_489 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_488; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_490 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_489; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_491 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_490; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_492 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_491; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_493 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_492; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_494 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_493; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_495 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_494; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_496 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_495; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_497 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_496; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_498 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_497; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_499 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_498; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_500 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_499; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_501 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_500; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_502 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_501; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_503 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_502; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_504 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_503; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_505 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_504; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_506 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_505; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_507 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_506; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_508 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_507; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_509 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_508; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_510 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_509; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_511 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_510; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_573 = 8'h3d == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_574 = 8'h3e == io_inputs_0[7:0] ? 7'ha : _GEN_573; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_575 = 8'h3f == io_inputs_0[7:0] ? 7'hf : _GEN_574; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_576 = 8'h40 == io_inputs_0[7:0] ? 7'h14 : _GEN_575; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_577 = 8'h41 == io_inputs_0[7:0] ? 7'h19 : _GEN_576; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_578 = 8'h42 == io_inputs_0[7:0] ? 7'h1e : _GEN_577; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_579 = 8'h43 == io_inputs_0[7:0] ? 7'h23 : _GEN_578; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_580 = 8'h44 == io_inputs_0[7:0] ? 7'h28 : _GEN_579; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_581 = 8'h45 == io_inputs_0[7:0] ? 7'h2d : _GEN_580; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_582 = 8'h46 == io_inputs_0[7:0] ? 7'h32 : _GEN_581; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_583 = 8'h47 == io_inputs_0[7:0] ? 7'h37 : _GEN_582; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_584 = 8'h48 == io_inputs_0[7:0] ? 7'h3c : _GEN_583; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_585 = 8'h49 == io_inputs_0[7:0] ? 7'h41 : _GEN_584; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_586 = 8'h4a == io_inputs_0[7:0] ? 7'h46 : _GEN_585; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_587 = 8'h4b == io_inputs_0[7:0] ? 7'h4b : _GEN_586; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_588 = 8'h4c == io_inputs_0[7:0] ? 7'h50 : _GEN_587; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_589 = 8'h4d == io_inputs_0[7:0] ? 7'h55 : _GEN_588; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_590 = 8'h4e == io_inputs_0[7:0] ? 7'h5a : _GEN_589; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_591 = 8'h4f == io_inputs_0[7:0] ? 7'h5f : _GEN_590; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_592 = 8'h50 == io_inputs_0[7:0] ? 7'h64 : _GEN_591; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_593 = 8'h51 == io_inputs_0[7:0] ? 7'h64 : _GEN_592; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_594 = 8'h52 == io_inputs_0[7:0] ? 7'h64 : _GEN_593; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_595 = 8'h53 == io_inputs_0[7:0] ? 7'h64 : _GEN_594; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_596 = 8'h54 == io_inputs_0[7:0] ? 7'h64 : _GEN_595; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_597 = 8'h55 == io_inputs_0[7:0] ? 7'h64 : _GEN_596; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_598 = 8'h56 == io_inputs_0[7:0] ? 7'h64 : _GEN_597; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_599 = 8'h57 == io_inputs_0[7:0] ? 7'h64 : _GEN_598; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_600 = 8'h58 == io_inputs_0[7:0] ? 7'h64 : _GEN_599; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_601 = 8'h59 == io_inputs_0[7:0] ? 7'h64 : _GEN_600; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_602 = 8'h5a == io_inputs_0[7:0] ? 7'h64 : _GEN_601; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_603 = 8'h5b == io_inputs_0[7:0] ? 7'h64 : _GEN_602; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_604 = 8'h5c == io_inputs_0[7:0] ? 7'h64 : _GEN_603; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_605 = 8'h5d == io_inputs_0[7:0] ? 7'h64 : _GEN_604; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_606 = 8'h5e == io_inputs_0[7:0] ? 7'h64 : _GEN_605; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_607 = 8'h5f == io_inputs_0[7:0] ? 7'h64 : _GEN_606; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_608 = 8'h60 == io_inputs_0[7:0] ? 7'h64 : _GEN_607; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_609 = 8'h61 == io_inputs_0[7:0] ? 7'h64 : _GEN_608; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_610 = 8'h62 == io_inputs_0[7:0] ? 7'h64 : _GEN_609; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_611 = 8'h63 == io_inputs_0[7:0] ? 7'h64 : _GEN_610; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_612 = 8'h64 == io_inputs_0[7:0] ? 7'h64 : _GEN_611; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_613 = 8'h65 == io_inputs_0[7:0] ? 7'h5f : _GEN_612; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_614 = 8'h66 == io_inputs_0[7:0] ? 7'h5a : _GEN_613; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_615 = 8'h67 == io_inputs_0[7:0] ? 7'h55 : _GEN_614; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_616 = 8'h68 == io_inputs_0[7:0] ? 7'h50 : _GEN_615; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_617 = 8'h69 == io_inputs_0[7:0] ? 7'h4b : _GEN_616; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_618 = 8'h6a == io_inputs_0[7:0] ? 7'h46 : _GEN_617; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_619 = 8'h6b == io_inputs_0[7:0] ? 7'h41 : _GEN_618; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_620 = 8'h6c == io_inputs_0[7:0] ? 7'h3c : _GEN_619; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_621 = 8'h6d == io_inputs_0[7:0] ? 7'h37 : _GEN_620; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_622 = 8'h6e == io_inputs_0[7:0] ? 7'h32 : _GEN_621; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_623 = 8'h6f == io_inputs_0[7:0] ? 7'h2d : _GEN_622; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_624 = 8'h70 == io_inputs_0[7:0] ? 7'h28 : _GEN_623; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_625 = 8'h71 == io_inputs_0[7:0] ? 7'h23 : _GEN_624; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_626 = 8'h72 == io_inputs_0[7:0] ? 7'h1e : _GEN_625; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_627 = 8'h73 == io_inputs_0[7:0] ? 7'h19 : _GEN_626; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_628 = 8'h74 == io_inputs_0[7:0] ? 7'h14 : _GEN_627; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_629 = 8'h75 == io_inputs_0[7:0] ? 7'hf : _GEN_628; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_630 = 8'h76 == io_inputs_0[7:0] ? 7'ha : _GEN_629; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_631 = 8'h77 == io_inputs_0[7:0] ? 7'h5 : _GEN_630; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_632 = 8'h78 == io_inputs_0[7:0] ? 7'h0 : _GEN_631; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_633 = 8'h79 == io_inputs_0[7:0] ? 7'h0 : _GEN_632; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_634 = 8'h7a == io_inputs_0[7:0] ? 7'h0 : _GEN_633; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_635 = 8'h7b == io_inputs_0[7:0] ? 7'h0 : _GEN_634; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_636 = 8'h7c == io_inputs_0[7:0] ? 7'h0 : _GEN_635; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_637 = 8'h7d == io_inputs_0[7:0] ? 7'h0 : _GEN_636; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_638 = 8'h7e == io_inputs_0[7:0] ? 7'h0 : _GEN_637; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_639 = 8'h7f == io_inputs_0[7:0] ? 7'h0 : _GEN_638; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_640 = 8'h80 == io_inputs_0[7:0] ? 7'h0 : _GEN_639; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_641 = 8'h81 == io_inputs_0[7:0] ? 7'h0 : _GEN_640; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_642 = 8'h82 == io_inputs_0[7:0] ? 7'h0 : _GEN_641; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_643 = 8'h83 == io_inputs_0[7:0] ? 7'h0 : _GEN_642; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_644 = 8'h84 == io_inputs_0[7:0] ? 7'h0 : _GEN_643; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_645 = 8'h85 == io_inputs_0[7:0] ? 7'h0 : _GEN_644; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_646 = 8'h86 == io_inputs_0[7:0] ? 7'h0 : _GEN_645; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_647 = 8'h87 == io_inputs_0[7:0] ? 7'h0 : _GEN_646; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_648 = 8'h88 == io_inputs_0[7:0] ? 7'h0 : _GEN_647; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_649 = 8'h89 == io_inputs_0[7:0] ? 7'h0 : _GEN_648; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_650 = 8'h8a == io_inputs_0[7:0] ? 7'h0 : _GEN_649; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_651 = 8'h8b == io_inputs_0[7:0] ? 7'h0 : _GEN_650; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_652 = 8'h8c == io_inputs_0[7:0] ? 7'h0 : _GEN_651; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_653 = 8'h8d == io_inputs_0[7:0] ? 7'h0 : _GEN_652; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_654 = 8'h8e == io_inputs_0[7:0] ? 7'h0 : _GEN_653; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_655 = 8'h8f == io_inputs_0[7:0] ? 7'h0 : _GEN_654; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_656 = 8'h90 == io_inputs_0[7:0] ? 7'h0 : _GEN_655; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_657 = 8'h91 == io_inputs_0[7:0] ? 7'h0 : _GEN_656; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_658 = 8'h92 == io_inputs_0[7:0] ? 7'h0 : _GEN_657; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_659 = 8'h93 == io_inputs_0[7:0] ? 7'h0 : _GEN_658; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_660 = 8'h94 == io_inputs_0[7:0] ? 7'h0 : _GEN_659; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_661 = 8'h95 == io_inputs_0[7:0] ? 7'h0 : _GEN_660; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_662 = 8'h96 == io_inputs_0[7:0] ? 7'h0 : _GEN_661; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_663 = 8'h97 == io_inputs_0[7:0] ? 7'h0 : _GEN_662; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_664 = 8'h98 == io_inputs_0[7:0] ? 7'h0 : _GEN_663; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_665 = 8'h99 == io_inputs_0[7:0] ? 7'h0 : _GEN_664; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_666 = 8'h9a == io_inputs_0[7:0] ? 7'h0 : _GEN_665; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_667 = 8'h9b == io_inputs_0[7:0] ? 7'h0 : _GEN_666; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_668 = 8'h9c == io_inputs_0[7:0] ? 7'h0 : _GEN_667; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_669 = 8'h9d == io_inputs_0[7:0] ? 7'h0 : _GEN_668; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_670 = 8'h9e == io_inputs_0[7:0] ? 7'h0 : _GEN_669; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_671 = 8'h9f == io_inputs_0[7:0] ? 7'h0 : _GEN_670; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_672 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_671; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_673 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_672; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_674 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_673; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_675 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_674; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_676 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_675; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_677 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_676; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_678 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_677; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_679 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_678; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_680 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_679; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_681 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_680; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_682 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_681; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_683 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_682; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_684 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_683; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_685 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_684; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_686 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_685; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_687 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_686; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_688 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_687; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_689 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_688; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_690 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_689; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_691 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_690; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_692 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_691; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_693 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_692; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_694 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_693; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_695 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_694; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_696 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_695; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_697 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_696; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_698 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_697; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_699 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_698; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_700 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_699; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_701 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_700; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_702 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_701; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_703 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_702; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_704 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_703; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_705 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_704; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_706 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_705; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_707 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_706; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_708 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_707; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_709 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_708; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_710 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_709; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_711 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_710; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_712 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_711; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_713 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_712; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_714 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_713; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_715 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_714; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_716 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_715; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_717 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_716; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_718 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_717; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_719 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_718; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_720 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_719; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_721 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_720; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_722 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_721; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_723 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_722; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_724 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_723; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_725 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_724; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_726 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_725; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_727 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_726; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_728 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_727; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_729 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_728; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_730 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_729; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_731 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_730; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_732 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_731; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_733 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_732; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_734 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_733; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_735 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_734; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_736 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_735; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_737 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_736; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_738 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_737; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_739 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_738; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_740 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_739; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_741 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_740; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_742 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_741; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_743 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_742; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_744 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_743; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_745 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_744; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_746 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_745; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_747 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_746; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_748 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_747; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_749 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_748; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_750 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_749; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_751 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_750; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_752 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_751; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_753 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_752; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_754 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_753; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_755 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_754; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_756 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_755; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_757 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_756; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_758 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_757; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_759 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_758; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_760 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_759; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_761 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_760; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_762 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_761; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_763 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_762; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_764 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_763; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_765 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_764; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_766 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_765; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_767 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_766; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_869 = 8'h65 == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_870 = 8'h66 == io_inputs_0[7:0] ? 7'ha : _GEN_869; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_871 = 8'h67 == io_inputs_0[7:0] ? 7'hf : _GEN_870; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_872 = 8'h68 == io_inputs_0[7:0] ? 7'h14 : _GEN_871; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_873 = 8'h69 == io_inputs_0[7:0] ? 7'h19 : _GEN_872; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_874 = 8'h6a == io_inputs_0[7:0] ? 7'h1e : _GEN_873; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_875 = 8'h6b == io_inputs_0[7:0] ? 7'h23 : _GEN_874; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_876 = 8'h6c == io_inputs_0[7:0] ? 7'h28 : _GEN_875; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_877 = 8'h6d == io_inputs_0[7:0] ? 7'h2d : _GEN_876; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_878 = 8'h6e == io_inputs_0[7:0] ? 7'h32 : _GEN_877; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_879 = 8'h6f == io_inputs_0[7:0] ? 7'h37 : _GEN_878; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_880 = 8'h70 == io_inputs_0[7:0] ? 7'h3c : _GEN_879; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_881 = 8'h71 == io_inputs_0[7:0] ? 7'h41 : _GEN_880; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_882 = 8'h72 == io_inputs_0[7:0] ? 7'h46 : _GEN_881; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_883 = 8'h73 == io_inputs_0[7:0] ? 7'h4b : _GEN_882; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_884 = 8'h74 == io_inputs_0[7:0] ? 7'h50 : _GEN_883; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_885 = 8'h75 == io_inputs_0[7:0] ? 7'h55 : _GEN_884; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_886 = 8'h76 == io_inputs_0[7:0] ? 7'h5a : _GEN_885; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_887 = 8'h77 == io_inputs_0[7:0] ? 7'h5f : _GEN_886; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_888 = 8'h78 == io_inputs_0[7:0] ? 7'h64 : _GEN_887; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_889 = 8'h79 == io_inputs_0[7:0] ? 7'h64 : _GEN_888; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_890 = 8'h7a == io_inputs_0[7:0] ? 7'h64 : _GEN_889; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_891 = 8'h7b == io_inputs_0[7:0] ? 7'h64 : _GEN_890; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_892 = 8'h7c == io_inputs_0[7:0] ? 7'h64 : _GEN_891; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_893 = 8'h7d == io_inputs_0[7:0] ? 7'h64 : _GEN_892; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_894 = 8'h7e == io_inputs_0[7:0] ? 7'h64 : _GEN_893; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_895 = 8'h7f == io_inputs_0[7:0] ? 7'h64 : _GEN_894; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_896 = 8'h80 == io_inputs_0[7:0] ? 7'h64 : _GEN_895; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_897 = 8'h81 == io_inputs_0[7:0] ? 7'h64 : _GEN_896; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_898 = 8'h82 == io_inputs_0[7:0] ? 7'h64 : _GEN_897; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_899 = 8'h83 == io_inputs_0[7:0] ? 7'h64 : _GEN_898; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_900 = 8'h84 == io_inputs_0[7:0] ? 7'h64 : _GEN_899; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_901 = 8'h85 == io_inputs_0[7:0] ? 7'h64 : _GEN_900; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_902 = 8'h86 == io_inputs_0[7:0] ? 7'h64 : _GEN_901; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_903 = 8'h87 == io_inputs_0[7:0] ? 7'h64 : _GEN_902; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_904 = 8'h88 == io_inputs_0[7:0] ? 7'h64 : _GEN_903; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_905 = 8'h89 == io_inputs_0[7:0] ? 7'h64 : _GEN_904; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_906 = 8'h8a == io_inputs_0[7:0] ? 7'h64 : _GEN_905; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_907 = 8'h8b == io_inputs_0[7:0] ? 7'h64 : _GEN_906; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_908 = 8'h8c == io_inputs_0[7:0] ? 7'h64 : _GEN_907; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_909 = 8'h8d == io_inputs_0[7:0] ? 7'h5f : _GEN_908; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_910 = 8'h8e == io_inputs_0[7:0] ? 7'h5a : _GEN_909; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_911 = 8'h8f == io_inputs_0[7:0] ? 7'h55 : _GEN_910; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_912 = 8'h90 == io_inputs_0[7:0] ? 7'h50 : _GEN_911; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_913 = 8'h91 == io_inputs_0[7:0] ? 7'h4b : _GEN_912; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_914 = 8'h92 == io_inputs_0[7:0] ? 7'h46 : _GEN_913; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_915 = 8'h93 == io_inputs_0[7:0] ? 7'h41 : _GEN_914; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_916 = 8'h94 == io_inputs_0[7:0] ? 7'h3c : _GEN_915; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_917 = 8'h95 == io_inputs_0[7:0] ? 7'h37 : _GEN_916; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_918 = 8'h96 == io_inputs_0[7:0] ? 7'h32 : _GEN_917; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_919 = 8'h97 == io_inputs_0[7:0] ? 7'h2d : _GEN_918; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_920 = 8'h98 == io_inputs_0[7:0] ? 7'h28 : _GEN_919; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_921 = 8'h99 == io_inputs_0[7:0] ? 7'h23 : _GEN_920; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_922 = 8'h9a == io_inputs_0[7:0] ? 7'h1e : _GEN_921; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_923 = 8'h9b == io_inputs_0[7:0] ? 7'h19 : _GEN_922; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_924 = 8'h9c == io_inputs_0[7:0] ? 7'h14 : _GEN_923; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_925 = 8'h9d == io_inputs_0[7:0] ? 7'hf : _GEN_924; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_926 = 8'h9e == io_inputs_0[7:0] ? 7'ha : _GEN_925; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_927 = 8'h9f == io_inputs_0[7:0] ? 7'h5 : _GEN_926; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_928 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_927; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_929 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_928; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_930 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_929; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_931 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_930; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_932 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_931; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_933 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_932; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_934 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_933; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_935 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_934; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_936 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_935; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_937 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_936; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_938 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_937; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_939 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_938; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_940 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_939; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_941 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_940; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_942 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_941; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_943 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_942; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_944 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_943; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_945 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_944; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_946 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_945; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_947 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_946; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_948 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_947; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_949 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_948; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_950 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_949; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_951 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_950; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_952 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_951; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_953 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_952; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_954 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_953; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_955 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_954; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_956 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_955; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_957 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_956; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_958 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_957; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_959 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_958; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_960 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_959; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_961 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_960; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_962 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_961; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_963 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_962; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_964 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_963; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_965 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_964; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_966 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_965; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_967 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_966; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_968 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_967; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_969 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_968; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_970 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_969; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_971 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_970; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_972 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_971; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_973 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_972; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_974 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_973; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_975 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_974; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_976 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_975; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_977 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_976; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_978 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_977; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_979 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_978; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_980 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_979; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_981 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_980; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_982 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_981; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_983 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_982; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_984 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_983; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_985 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_984; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_986 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_985; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_987 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_986; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_988 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_987; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_989 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_988; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_990 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_989; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_991 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_990; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_992 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_991; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_993 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_992; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_994 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_993; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_995 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_994; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_996 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_995; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_997 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_996; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_998 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_997; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_999 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_998; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1000 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_999; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1001 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_1000; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1002 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_1001; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1003 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_1002; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1004 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_1003; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1005 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_1004; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1006 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_1005; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1007 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_1006; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1008 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_1007; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1009 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_1008; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1010 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_1009; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1011 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_1010; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1012 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_1011; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1013 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_1012; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1014 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_1013; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1015 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_1014; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1016 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_1015; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1017 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_1016; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1018 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_1017; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1019 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_1018; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1020 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_1019; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1021 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_1020; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1022 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_1021; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1023 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_1022; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1165 = 8'h8d == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1166 = 8'h8e == io_inputs_0[7:0] ? 7'ha : _GEN_1165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1167 = 8'h8f == io_inputs_0[7:0] ? 7'hf : _GEN_1166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1168 = 8'h90 == io_inputs_0[7:0] ? 7'h14 : _GEN_1167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1169 = 8'h91 == io_inputs_0[7:0] ? 7'h19 : _GEN_1168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1170 = 8'h92 == io_inputs_0[7:0] ? 7'h1e : _GEN_1169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1171 = 8'h93 == io_inputs_0[7:0] ? 7'h23 : _GEN_1170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1172 = 8'h94 == io_inputs_0[7:0] ? 7'h28 : _GEN_1171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1173 = 8'h95 == io_inputs_0[7:0] ? 7'h2d : _GEN_1172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1174 = 8'h96 == io_inputs_0[7:0] ? 7'h32 : _GEN_1173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1175 = 8'h97 == io_inputs_0[7:0] ? 7'h37 : _GEN_1174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1176 = 8'h98 == io_inputs_0[7:0] ? 7'h3c : _GEN_1175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1177 = 8'h99 == io_inputs_0[7:0] ? 7'h41 : _GEN_1176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1178 = 8'h9a == io_inputs_0[7:0] ? 7'h46 : _GEN_1177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1179 = 8'h9b == io_inputs_0[7:0] ? 7'h4b : _GEN_1178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1180 = 8'h9c == io_inputs_0[7:0] ? 7'h50 : _GEN_1179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1181 = 8'h9d == io_inputs_0[7:0] ? 7'h55 : _GEN_1180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1182 = 8'h9e == io_inputs_0[7:0] ? 7'h5a : _GEN_1181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1183 = 8'h9f == io_inputs_0[7:0] ? 7'h5f : _GEN_1182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1184 = 8'ha0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1185 = 8'ha1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1186 = 8'ha2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1187 = 8'ha3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1188 = 8'ha4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1189 = 8'ha5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1190 = 8'ha6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1191 = 8'ha7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1192 = 8'ha8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1193 = 8'ha9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1194 = 8'haa == io_inputs_0[7:0] ? 7'h64 : _GEN_1193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1195 = 8'hab == io_inputs_0[7:0] ? 7'h64 : _GEN_1194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1196 = 8'hac == io_inputs_0[7:0] ? 7'h64 : _GEN_1195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1197 = 8'had == io_inputs_0[7:0] ? 7'h64 : _GEN_1196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1198 = 8'hae == io_inputs_0[7:0] ? 7'h64 : _GEN_1197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1199 = 8'haf == io_inputs_0[7:0] ? 7'h64 : _GEN_1198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1200 = 8'hb0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1201 = 8'hb1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1202 = 8'hb2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1203 = 8'hb3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1204 = 8'hb4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1205 = 8'hb5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1206 = 8'hb6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1207 = 8'hb7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1208 = 8'hb8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1209 = 8'hb9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1210 = 8'hba == io_inputs_0[7:0] ? 7'h64 : _GEN_1209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1211 = 8'hbb == io_inputs_0[7:0] ? 7'h64 : _GEN_1210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1212 = 8'hbc == io_inputs_0[7:0] ? 7'h64 : _GEN_1211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1213 = 8'hbd == io_inputs_0[7:0] ? 7'h64 : _GEN_1212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1214 = 8'hbe == io_inputs_0[7:0] ? 7'h64 : _GEN_1213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1215 = 8'hbf == io_inputs_0[7:0] ? 7'h64 : _GEN_1214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1216 = 8'hc0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1217 = 8'hc1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1218 = 8'hc2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1219 = 8'hc3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1220 = 8'hc4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1221 = 8'hc5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1222 = 8'hc6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1223 = 8'hc7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1224 = 8'hc8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1225 = 8'hc9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1226 = 8'hca == io_inputs_0[7:0] ? 7'h64 : _GEN_1225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1227 = 8'hcb == io_inputs_0[7:0] ? 7'h64 : _GEN_1226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1228 = 8'hcc == io_inputs_0[7:0] ? 7'h64 : _GEN_1227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1229 = 8'hcd == io_inputs_0[7:0] ? 7'h64 : _GEN_1228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1230 = 8'hce == io_inputs_0[7:0] ? 7'h64 : _GEN_1229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1231 = 8'hcf == io_inputs_0[7:0] ? 7'h64 : _GEN_1230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1232 = 8'hd0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1233 = 8'hd1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1234 = 8'hd2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1235 = 8'hd3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1236 = 8'hd4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1237 = 8'hd5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1238 = 8'hd6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1239 = 8'hd7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1240 = 8'hd8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1241 = 8'hd9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1242 = 8'hda == io_inputs_0[7:0] ? 7'h64 : _GEN_1241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1243 = 8'hdb == io_inputs_0[7:0] ? 7'h64 : _GEN_1242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1244 = 8'hdc == io_inputs_0[7:0] ? 7'h64 : _GEN_1243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1245 = 8'hdd == io_inputs_0[7:0] ? 7'h64 : _GEN_1244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1246 = 8'hde == io_inputs_0[7:0] ? 7'h64 : _GEN_1245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1247 = 8'hdf == io_inputs_0[7:0] ? 7'h64 : _GEN_1246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1248 = 8'he0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1249 = 8'he1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1250 = 8'he2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1251 = 8'he3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1252 = 8'he4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1253 = 8'he5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1254 = 8'he6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1255 = 8'he7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1256 = 8'he8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1255; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1257 = 8'he9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1256; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1258 = 8'hea == io_inputs_0[7:0] ? 7'h64 : _GEN_1257; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1259 = 8'heb == io_inputs_0[7:0] ? 7'h64 : _GEN_1258; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1260 = 8'hec == io_inputs_0[7:0] ? 7'h64 : _GEN_1259; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1261 = 8'hed == io_inputs_0[7:0] ? 7'h64 : _GEN_1260; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1262 = 8'hee == io_inputs_0[7:0] ? 7'h64 : _GEN_1261; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1263 = 8'hef == io_inputs_0[7:0] ? 7'h64 : _GEN_1262; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1264 = 8'hf0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1263; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1265 = 8'hf1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1264; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1266 = 8'hf2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1265; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1267 = 8'hf3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1266; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1268 = 8'hf4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1267; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1269 = 8'hf5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1268; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1270 = 8'hf6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1269; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1271 = 8'hf7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1270; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1272 = 8'hf8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1271; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1273 = 8'hf9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1272; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1274 = 8'hfa == io_inputs_0[7:0] ? 7'h64 : _GEN_1273; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1275 = 8'hfb == io_inputs_0[7:0] ? 7'h64 : _GEN_1274; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1276 = 8'hfc == io_inputs_0[7:0] ? 7'h64 : _GEN_1275; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1277 = 8'hfd == io_inputs_0[7:0] ? 7'h64 : _GEN_1276; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1278 = 8'hfe == io_inputs_0[7:0] ? 7'h64 : _GEN_1277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1279 = 8'hff == io_inputs_0[7:0] ? 7'h64 : _GEN_1278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1331 = 10'h33 == io_inputs_1 ? 7'h63 : 7'h64; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1332 = 10'h34 == io_inputs_1 ? 7'h62 : _GEN_1331; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1333 = 10'h35 == io_inputs_1 ? 7'h61 : _GEN_1332; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1334 = 10'h36 == io_inputs_1 ? 7'h60 : _GEN_1333; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1335 = 10'h37 == io_inputs_1 ? 7'h5f : _GEN_1334; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1336 = 10'h38 == io_inputs_1 ? 7'h5e : _GEN_1335; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1337 = 10'h39 == io_inputs_1 ? 7'h5d : _GEN_1336; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1338 = 10'h3a == io_inputs_1 ? 7'h5c : _GEN_1337; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1339 = 10'h3b == io_inputs_1 ? 7'h5b : _GEN_1338; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1340 = 10'h3c == io_inputs_1 ? 7'h5a : _GEN_1339; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1341 = 10'h3d == io_inputs_1 ? 7'h59 : _GEN_1340; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1342 = 10'h3e == io_inputs_1 ? 7'h58 : _GEN_1341; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1343 = 10'h3f == io_inputs_1 ? 7'h57 : _GEN_1342; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1344 = 10'h40 == io_inputs_1 ? 7'h56 : _GEN_1343; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1345 = 10'h41 == io_inputs_1 ? 7'h55 : _GEN_1344; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1346 = 10'h42 == io_inputs_1 ? 7'h54 : _GEN_1345; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1347 = 10'h43 == io_inputs_1 ? 7'h53 : _GEN_1346; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1348 = 10'h44 == io_inputs_1 ? 7'h52 : _GEN_1347; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1349 = 10'h45 == io_inputs_1 ? 7'h51 : _GEN_1348; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1350 = 10'h46 == io_inputs_1 ? 7'h50 : _GEN_1349; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1351 = 10'h47 == io_inputs_1 ? 7'h4f : _GEN_1350; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1352 = 10'h48 == io_inputs_1 ? 7'h4e : _GEN_1351; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1353 = 10'h49 == io_inputs_1 ? 7'h4d : _GEN_1352; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1354 = 10'h4a == io_inputs_1 ? 7'h4c : _GEN_1353; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1355 = 10'h4b == io_inputs_1 ? 7'h4b : _GEN_1354; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1356 = 10'h4c == io_inputs_1 ? 7'h4a : _GEN_1355; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1357 = 10'h4d == io_inputs_1 ? 7'h49 : _GEN_1356; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1358 = 10'h4e == io_inputs_1 ? 7'h48 : _GEN_1357; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1359 = 10'h4f == io_inputs_1 ? 7'h47 : _GEN_1358; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1360 = 10'h50 == io_inputs_1 ? 7'h46 : _GEN_1359; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1361 = 10'h51 == io_inputs_1 ? 7'h45 : _GEN_1360; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1362 = 10'h52 == io_inputs_1 ? 7'h44 : _GEN_1361; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1363 = 10'h53 == io_inputs_1 ? 7'h43 : _GEN_1362; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1364 = 10'h54 == io_inputs_1 ? 7'h42 : _GEN_1363; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1365 = 10'h55 == io_inputs_1 ? 7'h41 : _GEN_1364; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1366 = 10'h56 == io_inputs_1 ? 7'h40 : _GEN_1365; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1367 = 10'h57 == io_inputs_1 ? 7'h3f : _GEN_1366; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1368 = 10'h58 == io_inputs_1 ? 7'h3e : _GEN_1367; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1369 = 10'h59 == io_inputs_1 ? 7'h3d : _GEN_1368; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1370 = 10'h5a == io_inputs_1 ? 7'h3c : _GEN_1369; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1371 = 10'h5b == io_inputs_1 ? 7'h3b : _GEN_1370; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1372 = 10'h5c == io_inputs_1 ? 7'h3a : _GEN_1371; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1373 = 10'h5d == io_inputs_1 ? 7'h39 : _GEN_1372; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1374 = 10'h5e == io_inputs_1 ? 7'h38 : _GEN_1373; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1375 = 10'h5f == io_inputs_1 ? 7'h37 : _GEN_1374; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1376 = 10'h60 == io_inputs_1 ? 7'h36 : _GEN_1375; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1377 = 10'h61 == io_inputs_1 ? 7'h35 : _GEN_1376; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1378 = 10'h62 == io_inputs_1 ? 7'h34 : _GEN_1377; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1379 = 10'h63 == io_inputs_1 ? 7'h33 : _GEN_1378; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1380 = 10'h64 == io_inputs_1 ? 7'h32 : _GEN_1379; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1381 = 10'h65 == io_inputs_1 ? 7'h31 : _GEN_1380; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1382 = 10'h66 == io_inputs_1 ? 7'h30 : _GEN_1381; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1383 = 10'h67 == io_inputs_1 ? 7'h2f : _GEN_1382; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1384 = 10'h68 == io_inputs_1 ? 7'h2e : _GEN_1383; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1385 = 10'h69 == io_inputs_1 ? 7'h2d : _GEN_1384; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1386 = 10'h6a == io_inputs_1 ? 7'h2c : _GEN_1385; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1387 = 10'h6b == io_inputs_1 ? 7'h2b : _GEN_1386; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1388 = 10'h6c == io_inputs_1 ? 7'h2a : _GEN_1387; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1389 = 10'h6d == io_inputs_1 ? 7'h29 : _GEN_1388; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1390 = 10'h6e == io_inputs_1 ? 7'h28 : _GEN_1389; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1391 = 10'h6f == io_inputs_1 ? 7'h27 : _GEN_1390; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1392 = 10'h70 == io_inputs_1 ? 7'h26 : _GEN_1391; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1393 = 10'h71 == io_inputs_1 ? 7'h25 : _GEN_1392; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1394 = 10'h72 == io_inputs_1 ? 7'h24 : _GEN_1393; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1395 = 10'h73 == io_inputs_1 ? 7'h23 : _GEN_1394; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1396 = 10'h74 == io_inputs_1 ? 7'h22 : _GEN_1395; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1397 = 10'h75 == io_inputs_1 ? 7'h21 : _GEN_1396; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1398 = 10'h76 == io_inputs_1 ? 7'h20 : _GEN_1397; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1399 = 10'h77 == io_inputs_1 ? 7'h1f : _GEN_1398; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1400 = 10'h78 == io_inputs_1 ? 7'h1e : _GEN_1399; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1401 = 10'h79 == io_inputs_1 ? 7'h1d : _GEN_1400; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1402 = 10'h7a == io_inputs_1 ? 7'h1c : _GEN_1401; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1403 = 10'h7b == io_inputs_1 ? 7'h1b : _GEN_1402; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1404 = 10'h7c == io_inputs_1 ? 7'h1a : _GEN_1403; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1405 = 10'h7d == io_inputs_1 ? 7'h19 : _GEN_1404; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1406 = 10'h7e == io_inputs_1 ? 7'h18 : _GEN_1405; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1407 = 10'h7f == io_inputs_1 ? 7'h17 : _GEN_1406; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1408 = 10'h80 == io_inputs_1 ? 7'h16 : _GEN_1407; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1409 = 10'h81 == io_inputs_1 ? 7'h15 : _GEN_1408; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1410 = 10'h82 == io_inputs_1 ? 7'h14 : _GEN_1409; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1411 = 10'h83 == io_inputs_1 ? 7'h13 : _GEN_1410; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1412 = 10'h84 == io_inputs_1 ? 7'h12 : _GEN_1411; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1413 = 10'h85 == io_inputs_1 ? 7'h11 : _GEN_1412; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1414 = 10'h86 == io_inputs_1 ? 7'h10 : _GEN_1413; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1415 = 10'h87 == io_inputs_1 ? 7'hf : _GEN_1414; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1416 = 10'h88 == io_inputs_1 ? 7'he : _GEN_1415; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1417 = 10'h89 == io_inputs_1 ? 7'hd : _GEN_1416; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1418 = 10'h8a == io_inputs_1 ? 7'hc : _GEN_1417; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1419 = 10'h8b == io_inputs_1 ? 7'hb : _GEN_1418; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1420 = 10'h8c == io_inputs_1 ? 7'ha : _GEN_1419; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1421 = 10'h8d == io_inputs_1 ? 7'h9 : _GEN_1420; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1422 = 10'h8e == io_inputs_1 ? 7'h8 : _GEN_1421; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1423 = 10'h8f == io_inputs_1 ? 7'h7 : _GEN_1422; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1424 = 10'h90 == io_inputs_1 ? 7'h6 : _GEN_1423; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1425 = 10'h91 == io_inputs_1 ? 7'h5 : _GEN_1424; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1426 = 10'h92 == io_inputs_1 ? 7'h4 : _GEN_1425; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1427 = 10'h93 == io_inputs_1 ? 7'h3 : _GEN_1426; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1428 = 10'h94 == io_inputs_1 ? 7'h2 : _GEN_1427; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1429 = 10'h95 == io_inputs_1 ? 7'h1 : _GEN_1428; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1430 = 10'h96 == io_inputs_1 ? 7'h0 : _GEN_1429; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1431 = 10'h97 == io_inputs_1 ? 7'h0 : _GEN_1430; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1432 = 10'h98 == io_inputs_1 ? 7'h0 : _GEN_1431; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1433 = 10'h99 == io_inputs_1 ? 7'h0 : _GEN_1432; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1434 = 10'h9a == io_inputs_1 ? 7'h0 : _GEN_1433; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1435 = 10'h9b == io_inputs_1 ? 7'h0 : _GEN_1434; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1436 = 10'h9c == io_inputs_1 ? 7'h0 : _GEN_1435; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1437 = 10'h9d == io_inputs_1 ? 7'h0 : _GEN_1436; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1438 = 10'h9e == io_inputs_1 ? 7'h0 : _GEN_1437; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1439 = 10'h9f == io_inputs_1 ? 7'h0 : _GEN_1438; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1440 = 10'ha0 == io_inputs_1 ? 7'h0 : _GEN_1439; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1441 = 10'ha1 == io_inputs_1 ? 7'h0 : _GEN_1440; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1442 = 10'ha2 == io_inputs_1 ? 7'h0 : _GEN_1441; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1443 = 10'ha3 == io_inputs_1 ? 7'h0 : _GEN_1442; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1444 = 10'ha4 == io_inputs_1 ? 7'h0 : _GEN_1443; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1445 = 10'ha5 == io_inputs_1 ? 7'h0 : _GEN_1444; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1446 = 10'ha6 == io_inputs_1 ? 7'h0 : _GEN_1445; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1447 = 10'ha7 == io_inputs_1 ? 7'h0 : _GEN_1446; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1448 = 10'ha8 == io_inputs_1 ? 7'h0 : _GEN_1447; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1449 = 10'ha9 == io_inputs_1 ? 7'h0 : _GEN_1448; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1450 = 10'haa == io_inputs_1 ? 7'h0 : _GEN_1449; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1451 = 10'hab == io_inputs_1 ? 7'h0 : _GEN_1450; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1452 = 10'hac == io_inputs_1 ? 7'h0 : _GEN_1451; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1453 = 10'had == io_inputs_1 ? 7'h0 : _GEN_1452; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1454 = 10'hae == io_inputs_1 ? 7'h0 : _GEN_1453; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1455 = 10'haf == io_inputs_1 ? 7'h0 : _GEN_1454; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1456 = 10'hb0 == io_inputs_1 ? 7'h0 : _GEN_1455; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1457 = 10'hb1 == io_inputs_1 ? 7'h0 : _GEN_1456; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1458 = 10'hb2 == io_inputs_1 ? 7'h0 : _GEN_1457; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1459 = 10'hb3 == io_inputs_1 ? 7'h0 : _GEN_1458; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1460 = 10'hb4 == io_inputs_1 ? 7'h0 : _GEN_1459; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1461 = 10'hb5 == io_inputs_1 ? 7'h0 : _GEN_1460; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1462 = 10'hb6 == io_inputs_1 ? 7'h0 : _GEN_1461; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1463 = 10'hb7 == io_inputs_1 ? 7'h0 : _GEN_1462; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1464 = 10'hb8 == io_inputs_1 ? 7'h0 : _GEN_1463; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1465 = 10'hb9 == io_inputs_1 ? 7'h0 : _GEN_1464; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1466 = 10'hba == io_inputs_1 ? 7'h0 : _GEN_1465; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1467 = 10'hbb == io_inputs_1 ? 7'h0 : _GEN_1466; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1468 = 10'hbc == io_inputs_1 ? 7'h0 : _GEN_1467; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1469 = 10'hbd == io_inputs_1 ? 7'h0 : _GEN_1468; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1470 = 10'hbe == io_inputs_1 ? 7'h0 : _GEN_1469; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1471 = 10'hbf == io_inputs_1 ? 7'h0 : _GEN_1470; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1472 = 10'hc0 == io_inputs_1 ? 7'h0 : _GEN_1471; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1473 = 10'hc1 == io_inputs_1 ? 7'h0 : _GEN_1472; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1474 = 10'hc2 == io_inputs_1 ? 7'h0 : _GEN_1473; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1475 = 10'hc3 == io_inputs_1 ? 7'h0 : _GEN_1474; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1476 = 10'hc4 == io_inputs_1 ? 7'h0 : _GEN_1475; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1477 = 10'hc5 == io_inputs_1 ? 7'h0 : _GEN_1476; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1478 = 10'hc6 == io_inputs_1 ? 7'h0 : _GEN_1477; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1479 = 10'hc7 == io_inputs_1 ? 7'h0 : _GEN_1478; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1480 = 10'hc8 == io_inputs_1 ? 7'h0 : _GEN_1479; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1481 = 10'hc9 == io_inputs_1 ? 7'h0 : _GEN_1480; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1482 = 10'hca == io_inputs_1 ? 7'h0 : _GEN_1481; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1483 = 10'hcb == io_inputs_1 ? 7'h0 : _GEN_1482; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1484 = 10'hcc == io_inputs_1 ? 7'h0 : _GEN_1483; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1485 = 10'hcd == io_inputs_1 ? 7'h0 : _GEN_1484; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1486 = 10'hce == io_inputs_1 ? 7'h0 : _GEN_1485; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1487 = 10'hcf == io_inputs_1 ? 7'h0 : _GEN_1486; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1488 = 10'hd0 == io_inputs_1 ? 7'h0 : _GEN_1487; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1489 = 10'hd1 == io_inputs_1 ? 7'h0 : _GEN_1488; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1490 = 10'hd2 == io_inputs_1 ? 7'h0 : _GEN_1489; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1491 = 10'hd3 == io_inputs_1 ? 7'h0 : _GEN_1490; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1492 = 10'hd4 == io_inputs_1 ? 7'h0 : _GEN_1491; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1493 = 10'hd5 == io_inputs_1 ? 7'h0 : _GEN_1492; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1494 = 10'hd6 == io_inputs_1 ? 7'h0 : _GEN_1493; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1495 = 10'hd7 == io_inputs_1 ? 7'h0 : _GEN_1494; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1496 = 10'hd8 == io_inputs_1 ? 7'h0 : _GEN_1495; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1497 = 10'hd9 == io_inputs_1 ? 7'h0 : _GEN_1496; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1498 = 10'hda == io_inputs_1 ? 7'h0 : _GEN_1497; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1499 = 10'hdb == io_inputs_1 ? 7'h0 : _GEN_1498; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1500 = 10'hdc == io_inputs_1 ? 7'h0 : _GEN_1499; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1501 = 10'hdd == io_inputs_1 ? 7'h0 : _GEN_1500; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1502 = 10'hde == io_inputs_1 ? 7'h0 : _GEN_1501; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1503 = 10'hdf == io_inputs_1 ? 7'h0 : _GEN_1502; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1504 = 10'he0 == io_inputs_1 ? 7'h0 : _GEN_1503; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1505 = 10'he1 == io_inputs_1 ? 7'h0 : _GEN_1504; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1506 = 10'he2 == io_inputs_1 ? 7'h0 : _GEN_1505; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1507 = 10'he3 == io_inputs_1 ? 7'h0 : _GEN_1506; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1508 = 10'he4 == io_inputs_1 ? 7'h0 : _GEN_1507; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1509 = 10'he5 == io_inputs_1 ? 7'h0 : _GEN_1508; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1510 = 10'he6 == io_inputs_1 ? 7'h0 : _GEN_1509; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1511 = 10'he7 == io_inputs_1 ? 7'h0 : _GEN_1510; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1512 = 10'he8 == io_inputs_1 ? 7'h0 : _GEN_1511; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1513 = 10'he9 == io_inputs_1 ? 7'h0 : _GEN_1512; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1514 = 10'hea == io_inputs_1 ? 7'h0 : _GEN_1513; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1515 = 10'heb == io_inputs_1 ? 7'h0 : _GEN_1514; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1516 = 10'hec == io_inputs_1 ? 7'h0 : _GEN_1515; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1517 = 10'hed == io_inputs_1 ? 7'h0 : _GEN_1516; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1518 = 10'hee == io_inputs_1 ? 7'h0 : _GEN_1517; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1519 = 10'hef == io_inputs_1 ? 7'h0 : _GEN_1518; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1520 = 10'hf0 == io_inputs_1 ? 7'h0 : _GEN_1519; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1521 = 10'hf1 == io_inputs_1 ? 7'h0 : _GEN_1520; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1522 = 10'hf2 == io_inputs_1 ? 7'h0 : _GEN_1521; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1523 = 10'hf3 == io_inputs_1 ? 7'h0 : _GEN_1522; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1524 = 10'hf4 == io_inputs_1 ? 7'h0 : _GEN_1523; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1525 = 10'hf5 == io_inputs_1 ? 7'h0 : _GEN_1524; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1526 = 10'hf6 == io_inputs_1 ? 7'h0 : _GEN_1525; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1527 = 10'hf7 == io_inputs_1 ? 7'h0 : _GEN_1526; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1528 = 10'hf8 == io_inputs_1 ? 7'h0 : _GEN_1527; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1529 = 10'hf9 == io_inputs_1 ? 7'h0 : _GEN_1528; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1530 = 10'hfa == io_inputs_1 ? 7'h0 : _GEN_1529; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1531 = 10'hfb == io_inputs_1 ? 7'h0 : _GEN_1530; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1532 = 10'hfc == io_inputs_1 ? 7'h0 : _GEN_1531; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1533 = 10'hfd == io_inputs_1 ? 7'h0 : _GEN_1532; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1534 = 10'hfe == io_inputs_1 ? 7'h0 : _GEN_1533; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1535 = 10'hff == io_inputs_1 ? 7'h0 : _GEN_1534; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1536 = 10'h100 == io_inputs_1 ? 7'h0 : _GEN_1535; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1537 = 10'h101 == io_inputs_1 ? 7'h0 : _GEN_1536; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1538 = 10'h102 == io_inputs_1 ? 7'h0 : _GEN_1537; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1539 = 10'h103 == io_inputs_1 ? 7'h0 : _GEN_1538; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1540 = 10'h104 == io_inputs_1 ? 7'h0 : _GEN_1539; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1541 = 10'h105 == io_inputs_1 ? 7'h0 : _GEN_1540; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1542 = 10'h106 == io_inputs_1 ? 7'h0 : _GEN_1541; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1543 = 10'h107 == io_inputs_1 ? 7'h0 : _GEN_1542; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1544 = 10'h108 == io_inputs_1 ? 7'h0 : _GEN_1543; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1545 = 10'h109 == io_inputs_1 ? 7'h0 : _GEN_1544; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1546 = 10'h10a == io_inputs_1 ? 7'h0 : _GEN_1545; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1547 = 10'h10b == io_inputs_1 ? 7'h0 : _GEN_1546; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1548 = 10'h10c == io_inputs_1 ? 7'h0 : _GEN_1547; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1549 = 10'h10d == io_inputs_1 ? 7'h0 : _GEN_1548; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1550 = 10'h10e == io_inputs_1 ? 7'h0 : _GEN_1549; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1551 = 10'h10f == io_inputs_1 ? 7'h0 : _GEN_1550; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1552 = 10'h110 == io_inputs_1 ? 7'h0 : _GEN_1551; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1553 = 10'h111 == io_inputs_1 ? 7'h0 : _GEN_1552; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1554 = 10'h112 == io_inputs_1 ? 7'h0 : _GEN_1553; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1555 = 10'h113 == io_inputs_1 ? 7'h0 : _GEN_1554; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1556 = 10'h114 == io_inputs_1 ? 7'h0 : _GEN_1555; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1557 = 10'h115 == io_inputs_1 ? 7'h0 : _GEN_1556; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1558 = 10'h116 == io_inputs_1 ? 7'h0 : _GEN_1557; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1559 = 10'h117 == io_inputs_1 ? 7'h0 : _GEN_1558; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1560 = 10'h118 == io_inputs_1 ? 7'h0 : _GEN_1559; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1561 = 10'h119 == io_inputs_1 ? 7'h0 : _GEN_1560; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1562 = 10'h11a == io_inputs_1 ? 7'h0 : _GEN_1561; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1563 = 10'h11b == io_inputs_1 ? 7'h0 : _GEN_1562; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1564 = 10'h11c == io_inputs_1 ? 7'h0 : _GEN_1563; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1565 = 10'h11d == io_inputs_1 ? 7'h0 : _GEN_1564; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1566 = 10'h11e == io_inputs_1 ? 7'h0 : _GEN_1565; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1567 = 10'h11f == io_inputs_1 ? 7'h0 : _GEN_1566; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1568 = 10'h120 == io_inputs_1 ? 7'h0 : _GEN_1567; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1569 = 10'h121 == io_inputs_1 ? 7'h0 : _GEN_1568; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1570 = 10'h122 == io_inputs_1 ? 7'h0 : _GEN_1569; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1571 = 10'h123 == io_inputs_1 ? 7'h0 : _GEN_1570; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1572 = 10'h124 == io_inputs_1 ? 7'h0 : _GEN_1571; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1573 = 10'h125 == io_inputs_1 ? 7'h0 : _GEN_1572; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1574 = 10'h126 == io_inputs_1 ? 7'h0 : _GEN_1573; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1575 = 10'h127 == io_inputs_1 ? 7'h0 : _GEN_1574; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1576 = 10'h128 == io_inputs_1 ? 7'h0 : _GEN_1575; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1577 = 10'h129 == io_inputs_1 ? 7'h0 : _GEN_1576; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1578 = 10'h12a == io_inputs_1 ? 7'h0 : _GEN_1577; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1579 = 10'h12b == io_inputs_1 ? 7'h0 : _GEN_1578; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1580 = 10'h12c == io_inputs_1 ? 7'h0 : _GEN_1579; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1581 = 10'h12d == io_inputs_1 ? 7'h0 : _GEN_1580; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1582 = 10'h12e == io_inputs_1 ? 7'h0 : _GEN_1581; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1583 = 10'h12f == io_inputs_1 ? 7'h0 : _GEN_1582; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1584 = 10'h130 == io_inputs_1 ? 7'h0 : _GEN_1583; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1585 = 10'h131 == io_inputs_1 ? 7'h0 : _GEN_1584; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1586 = 10'h132 == io_inputs_1 ? 7'h0 : _GEN_1585; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1587 = 10'h133 == io_inputs_1 ? 7'h0 : _GEN_1586; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1588 = 10'h134 == io_inputs_1 ? 7'h0 : _GEN_1587; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1589 = 10'h135 == io_inputs_1 ? 7'h0 : _GEN_1588; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1590 = 10'h136 == io_inputs_1 ? 7'h0 : _GEN_1589; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1591 = 10'h137 == io_inputs_1 ? 7'h0 : _GEN_1590; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1592 = 10'h138 == io_inputs_1 ? 7'h0 : _GEN_1591; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1593 = 10'h139 == io_inputs_1 ? 7'h0 : _GEN_1592; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1594 = 10'h13a == io_inputs_1 ? 7'h0 : _GEN_1593; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1595 = 10'h13b == io_inputs_1 ? 7'h0 : _GEN_1594; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1596 = 10'h13c == io_inputs_1 ? 7'h0 : _GEN_1595; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1597 = 10'h13d == io_inputs_1 ? 7'h0 : _GEN_1596; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1598 = 10'h13e == io_inputs_1 ? 7'h0 : _GEN_1597; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1599 = 10'h13f == io_inputs_1 ? 7'h0 : _GEN_1598; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1600 = 10'h140 == io_inputs_1 ? 7'h0 : _GEN_1599; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1601 = 10'h141 == io_inputs_1 ? 7'h0 : _GEN_1600; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1602 = 10'h142 == io_inputs_1 ? 7'h0 : _GEN_1601; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1603 = 10'h143 == io_inputs_1 ? 7'h0 : _GEN_1602; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1604 = 10'h144 == io_inputs_1 ? 7'h0 : _GEN_1603; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1605 = 10'h145 == io_inputs_1 ? 7'h0 : _GEN_1604; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1606 = 10'h146 == io_inputs_1 ? 7'h0 : _GEN_1605; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1607 = 10'h147 == io_inputs_1 ? 7'h0 : _GEN_1606; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1608 = 10'h148 == io_inputs_1 ? 7'h0 : _GEN_1607; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1609 = 10'h149 == io_inputs_1 ? 7'h0 : _GEN_1608; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1610 = 10'h14a == io_inputs_1 ? 7'h0 : _GEN_1609; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1611 = 10'h14b == io_inputs_1 ? 7'h0 : _GEN_1610; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1612 = 10'h14c == io_inputs_1 ? 7'h0 : _GEN_1611; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1613 = 10'h14d == io_inputs_1 ? 7'h0 : _GEN_1612; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1614 = 10'h14e == io_inputs_1 ? 7'h0 : _GEN_1613; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1615 = 10'h14f == io_inputs_1 ? 7'h0 : _GEN_1614; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1616 = 10'h150 == io_inputs_1 ? 7'h0 : _GEN_1615; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1617 = 10'h151 == io_inputs_1 ? 7'h0 : _GEN_1616; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1618 = 10'h152 == io_inputs_1 ? 7'h0 : _GEN_1617; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1619 = 10'h153 == io_inputs_1 ? 7'h0 : _GEN_1618; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1620 = 10'h154 == io_inputs_1 ? 7'h0 : _GEN_1619; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1621 = 10'h155 == io_inputs_1 ? 7'h0 : _GEN_1620; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1622 = 10'h156 == io_inputs_1 ? 7'h0 : _GEN_1621; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1623 = 10'h157 == io_inputs_1 ? 7'h0 : _GEN_1622; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1624 = 10'h158 == io_inputs_1 ? 7'h0 : _GEN_1623; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1625 = 10'h159 == io_inputs_1 ? 7'h0 : _GEN_1624; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1626 = 10'h15a == io_inputs_1 ? 7'h0 : _GEN_1625; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1627 = 10'h15b == io_inputs_1 ? 7'h0 : _GEN_1626; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1628 = 10'h15c == io_inputs_1 ? 7'h0 : _GEN_1627; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1629 = 10'h15d == io_inputs_1 ? 7'h0 : _GEN_1628; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1630 = 10'h15e == io_inputs_1 ? 7'h0 : _GEN_1629; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1631 = 10'h15f == io_inputs_1 ? 7'h0 : _GEN_1630; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1632 = 10'h160 == io_inputs_1 ? 7'h0 : _GEN_1631; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1633 = 10'h161 == io_inputs_1 ? 7'h0 : _GEN_1632; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1634 = 10'h162 == io_inputs_1 ? 7'h0 : _GEN_1633; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1635 = 10'h163 == io_inputs_1 ? 7'h0 : _GEN_1634; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1636 = 10'h164 == io_inputs_1 ? 7'h0 : _GEN_1635; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1637 = 10'h165 == io_inputs_1 ? 7'h0 : _GEN_1636; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1638 = 10'h166 == io_inputs_1 ? 7'h0 : _GEN_1637; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1639 = 10'h167 == io_inputs_1 ? 7'h0 : _GEN_1638; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1640 = 10'h168 == io_inputs_1 ? 7'h0 : _GEN_1639; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1641 = 10'h169 == io_inputs_1 ? 7'h0 : _GEN_1640; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1642 = 10'h16a == io_inputs_1 ? 7'h0 : _GEN_1641; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1643 = 10'h16b == io_inputs_1 ? 7'h0 : _GEN_1642; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1644 = 10'h16c == io_inputs_1 ? 7'h0 : _GEN_1643; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1645 = 10'h16d == io_inputs_1 ? 7'h0 : _GEN_1644; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1646 = 10'h16e == io_inputs_1 ? 7'h0 : _GEN_1645; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1647 = 10'h16f == io_inputs_1 ? 7'h0 : _GEN_1646; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1648 = 10'h170 == io_inputs_1 ? 7'h0 : _GEN_1647; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1649 = 10'h171 == io_inputs_1 ? 7'h0 : _GEN_1648; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1650 = 10'h172 == io_inputs_1 ? 7'h0 : _GEN_1649; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1651 = 10'h173 == io_inputs_1 ? 7'h0 : _GEN_1650; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1652 = 10'h174 == io_inputs_1 ? 7'h0 : _GEN_1651; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1653 = 10'h175 == io_inputs_1 ? 7'h0 : _GEN_1652; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1654 = 10'h176 == io_inputs_1 ? 7'h0 : _GEN_1653; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1655 = 10'h177 == io_inputs_1 ? 7'h0 : _GEN_1654; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1656 = 10'h178 == io_inputs_1 ? 7'h0 : _GEN_1655; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1657 = 10'h179 == io_inputs_1 ? 7'h0 : _GEN_1656; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1658 = 10'h17a == io_inputs_1 ? 7'h0 : _GEN_1657; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1659 = 10'h17b == io_inputs_1 ? 7'h0 : _GEN_1658; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1660 = 10'h17c == io_inputs_1 ? 7'h0 : _GEN_1659; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1661 = 10'h17d == io_inputs_1 ? 7'h0 : _GEN_1660; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1662 = 10'h17e == io_inputs_1 ? 7'h0 : _GEN_1661; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1663 = 10'h17f == io_inputs_1 ? 7'h0 : _GEN_1662; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1664 = 10'h180 == io_inputs_1 ? 7'h0 : _GEN_1663; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1665 = 10'h181 == io_inputs_1 ? 7'h0 : _GEN_1664; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1666 = 10'h182 == io_inputs_1 ? 7'h0 : _GEN_1665; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1667 = 10'h183 == io_inputs_1 ? 7'h0 : _GEN_1666; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1668 = 10'h184 == io_inputs_1 ? 7'h0 : _GEN_1667; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1669 = 10'h185 == io_inputs_1 ? 7'h0 : _GEN_1668; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1670 = 10'h186 == io_inputs_1 ? 7'h0 : _GEN_1669; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1671 = 10'h187 == io_inputs_1 ? 7'h0 : _GEN_1670; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1672 = 10'h188 == io_inputs_1 ? 7'h0 : _GEN_1671; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1673 = 10'h189 == io_inputs_1 ? 7'h0 : _GEN_1672; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1674 = 10'h18a == io_inputs_1 ? 7'h0 : _GEN_1673; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1675 = 10'h18b == io_inputs_1 ? 7'h0 : _GEN_1674; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1676 = 10'h18c == io_inputs_1 ? 7'h0 : _GEN_1675; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1677 = 10'h18d == io_inputs_1 ? 7'h0 : _GEN_1676; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1678 = 10'h18e == io_inputs_1 ? 7'h0 : _GEN_1677; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1679 = 10'h18f == io_inputs_1 ? 7'h0 : _GEN_1678; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1680 = 10'h190 == io_inputs_1 ? 7'h0 : _GEN_1679; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1681 = 10'h191 == io_inputs_1 ? 7'h0 : _GEN_1680; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1682 = 10'h192 == io_inputs_1 ? 7'h0 : _GEN_1681; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1683 = 10'h193 == io_inputs_1 ? 7'h0 : _GEN_1682; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1684 = 10'h194 == io_inputs_1 ? 7'h0 : _GEN_1683; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1685 = 10'h195 == io_inputs_1 ? 7'h0 : _GEN_1684; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1686 = 10'h196 == io_inputs_1 ? 7'h0 : _GEN_1685; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1687 = 10'h197 == io_inputs_1 ? 7'h0 : _GEN_1686; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1688 = 10'h198 == io_inputs_1 ? 7'h0 : _GEN_1687; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1689 = 10'h199 == io_inputs_1 ? 7'h0 : _GEN_1688; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1690 = 10'h19a == io_inputs_1 ? 7'h0 : _GEN_1689; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1691 = 10'h19b == io_inputs_1 ? 7'h0 : _GEN_1690; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1692 = 10'h19c == io_inputs_1 ? 7'h0 : _GEN_1691; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1693 = 10'h19d == io_inputs_1 ? 7'h0 : _GEN_1692; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1694 = 10'h19e == io_inputs_1 ? 7'h0 : _GEN_1693; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1695 = 10'h19f == io_inputs_1 ? 7'h0 : _GEN_1694; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1696 = 10'h1a0 == io_inputs_1 ? 7'h0 : _GEN_1695; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1697 = 10'h1a1 == io_inputs_1 ? 7'h0 : _GEN_1696; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1698 = 10'h1a2 == io_inputs_1 ? 7'h0 : _GEN_1697; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1699 = 10'h1a3 == io_inputs_1 ? 7'h0 : _GEN_1698; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1700 = 10'h1a4 == io_inputs_1 ? 7'h0 : _GEN_1699; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1701 = 10'h1a5 == io_inputs_1 ? 7'h0 : _GEN_1700; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1702 = 10'h1a6 == io_inputs_1 ? 7'h0 : _GEN_1701; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1703 = 10'h1a7 == io_inputs_1 ? 7'h0 : _GEN_1702; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1704 = 10'h1a8 == io_inputs_1 ? 7'h0 : _GEN_1703; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1705 = 10'h1a9 == io_inputs_1 ? 7'h0 : _GEN_1704; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1706 = 10'h1aa == io_inputs_1 ? 7'h0 : _GEN_1705; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1707 = 10'h1ab == io_inputs_1 ? 7'h0 : _GEN_1706; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1708 = 10'h1ac == io_inputs_1 ? 7'h0 : _GEN_1707; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1709 = 10'h1ad == io_inputs_1 ? 7'h0 : _GEN_1708; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1710 = 10'h1ae == io_inputs_1 ? 7'h0 : _GEN_1709; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1711 = 10'h1af == io_inputs_1 ? 7'h0 : _GEN_1710; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1712 = 10'h1b0 == io_inputs_1 ? 7'h0 : _GEN_1711; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1713 = 10'h1b1 == io_inputs_1 ? 7'h0 : _GEN_1712; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1714 = 10'h1b2 == io_inputs_1 ? 7'h0 : _GEN_1713; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1715 = 10'h1b3 == io_inputs_1 ? 7'h0 : _GEN_1714; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1716 = 10'h1b4 == io_inputs_1 ? 7'h0 : _GEN_1715; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1717 = 10'h1b5 == io_inputs_1 ? 7'h0 : _GEN_1716; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1718 = 10'h1b6 == io_inputs_1 ? 7'h0 : _GEN_1717; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1719 = 10'h1b7 == io_inputs_1 ? 7'h0 : _GEN_1718; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1720 = 10'h1b8 == io_inputs_1 ? 7'h0 : _GEN_1719; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1721 = 10'h1b9 == io_inputs_1 ? 7'h0 : _GEN_1720; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1722 = 10'h1ba == io_inputs_1 ? 7'h0 : _GEN_1721; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1723 = 10'h1bb == io_inputs_1 ? 7'h0 : _GEN_1722; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1724 = 10'h1bc == io_inputs_1 ? 7'h0 : _GEN_1723; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1725 = 10'h1bd == io_inputs_1 ? 7'h0 : _GEN_1724; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1726 = 10'h1be == io_inputs_1 ? 7'h0 : _GEN_1725; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1727 = 10'h1bf == io_inputs_1 ? 7'h0 : _GEN_1726; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1728 = 10'h1c0 == io_inputs_1 ? 7'h0 : _GEN_1727; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1729 = 10'h1c1 == io_inputs_1 ? 7'h0 : _GEN_1728; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1730 = 10'h1c2 == io_inputs_1 ? 7'h0 : _GEN_1729; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1731 = 10'h1c3 == io_inputs_1 ? 7'h0 : _GEN_1730; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1732 = 10'h1c4 == io_inputs_1 ? 7'h0 : _GEN_1731; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1733 = 10'h1c5 == io_inputs_1 ? 7'h0 : _GEN_1732; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1734 = 10'h1c6 == io_inputs_1 ? 7'h0 : _GEN_1733; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1735 = 10'h1c7 == io_inputs_1 ? 7'h0 : _GEN_1734; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1736 = 10'h1c8 == io_inputs_1 ? 7'h0 : _GEN_1735; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1737 = 10'h1c9 == io_inputs_1 ? 7'h0 : _GEN_1736; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1738 = 10'h1ca == io_inputs_1 ? 7'h0 : _GEN_1737; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1739 = 10'h1cb == io_inputs_1 ? 7'h0 : _GEN_1738; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1740 = 10'h1cc == io_inputs_1 ? 7'h0 : _GEN_1739; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1741 = 10'h1cd == io_inputs_1 ? 7'h0 : _GEN_1740; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1742 = 10'h1ce == io_inputs_1 ? 7'h0 : _GEN_1741; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1743 = 10'h1cf == io_inputs_1 ? 7'h0 : _GEN_1742; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1744 = 10'h1d0 == io_inputs_1 ? 7'h0 : _GEN_1743; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1745 = 10'h1d1 == io_inputs_1 ? 7'h0 : _GEN_1744; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1746 = 10'h1d2 == io_inputs_1 ? 7'h0 : _GEN_1745; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1747 = 10'h1d3 == io_inputs_1 ? 7'h0 : _GEN_1746; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1748 = 10'h1d4 == io_inputs_1 ? 7'h0 : _GEN_1747; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1749 = 10'h1d5 == io_inputs_1 ? 7'h0 : _GEN_1748; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1750 = 10'h1d6 == io_inputs_1 ? 7'h0 : _GEN_1749; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1751 = 10'h1d7 == io_inputs_1 ? 7'h0 : _GEN_1750; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1752 = 10'h1d8 == io_inputs_1 ? 7'h0 : _GEN_1751; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1753 = 10'h1d9 == io_inputs_1 ? 7'h0 : _GEN_1752; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1754 = 10'h1da == io_inputs_1 ? 7'h0 : _GEN_1753; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1755 = 10'h1db == io_inputs_1 ? 7'h0 : _GEN_1754; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1756 = 10'h1dc == io_inputs_1 ? 7'h0 : _GEN_1755; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1757 = 10'h1dd == io_inputs_1 ? 7'h0 : _GEN_1756; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1758 = 10'h1de == io_inputs_1 ? 7'h0 : _GEN_1757; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1759 = 10'h1df == io_inputs_1 ? 7'h0 : _GEN_1758; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1760 = 10'h1e0 == io_inputs_1 ? 7'h0 : _GEN_1759; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1761 = 10'h1e1 == io_inputs_1 ? 7'h0 : _GEN_1760; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1762 = 10'h1e2 == io_inputs_1 ? 7'h0 : _GEN_1761; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1763 = 10'h1e3 == io_inputs_1 ? 7'h0 : _GEN_1762; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1764 = 10'h1e4 == io_inputs_1 ? 7'h0 : _GEN_1763; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1765 = 10'h1e5 == io_inputs_1 ? 7'h0 : _GEN_1764; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1766 = 10'h1e6 == io_inputs_1 ? 7'h0 : _GEN_1765; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1767 = 10'h1e7 == io_inputs_1 ? 7'h0 : _GEN_1766; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1768 = 10'h1e8 == io_inputs_1 ? 7'h0 : _GEN_1767; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1769 = 10'h1e9 == io_inputs_1 ? 7'h0 : _GEN_1768; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1770 = 10'h1ea == io_inputs_1 ? 7'h0 : _GEN_1769; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1771 = 10'h1eb == io_inputs_1 ? 7'h0 : _GEN_1770; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1772 = 10'h1ec == io_inputs_1 ? 7'h0 : _GEN_1771; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1773 = 10'h1ed == io_inputs_1 ? 7'h0 : _GEN_1772; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1774 = 10'h1ee == io_inputs_1 ? 7'h0 : _GEN_1773; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1775 = 10'h1ef == io_inputs_1 ? 7'h0 : _GEN_1774; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1776 = 10'h1f0 == io_inputs_1 ? 7'h0 : _GEN_1775; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1777 = 10'h1f1 == io_inputs_1 ? 7'h0 : _GEN_1776; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1778 = 10'h1f2 == io_inputs_1 ? 7'h0 : _GEN_1777; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1779 = 10'h1f3 == io_inputs_1 ? 7'h0 : _GEN_1778; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1780 = 10'h1f4 == io_inputs_1 ? 7'h0 : _GEN_1779; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1781 = 10'h1f5 == io_inputs_1 ? 7'h0 : _GEN_1780; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1782 = 10'h1f6 == io_inputs_1 ? 7'h0 : _GEN_1781; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1783 = 10'h1f7 == io_inputs_1 ? 7'h0 : _GEN_1782; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1784 = 10'h1f8 == io_inputs_1 ? 7'h0 : _GEN_1783; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1785 = 10'h1f9 == io_inputs_1 ? 7'h0 : _GEN_1784; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1786 = 10'h1fa == io_inputs_1 ? 7'h0 : _GEN_1785; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1787 = 10'h1fb == io_inputs_1 ? 7'h0 : _GEN_1786; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1788 = 10'h1fc == io_inputs_1 ? 7'h0 : _GEN_1787; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1789 = 10'h1fd == io_inputs_1 ? 7'h0 : _GEN_1788; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1790 = 10'h1fe == io_inputs_1 ? 7'h0 : _GEN_1789; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1791 = 10'h1ff == io_inputs_1 ? 7'h0 : _GEN_1790; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1792 = 10'h200 == io_inputs_1 ? 7'h0 : _GEN_1791; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1793 = 10'h201 == io_inputs_1 ? 7'h0 : _GEN_1792; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1794 = 10'h202 == io_inputs_1 ? 7'h0 : _GEN_1793; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1795 = 10'h203 == io_inputs_1 ? 7'h0 : _GEN_1794; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1796 = 10'h204 == io_inputs_1 ? 7'h0 : _GEN_1795; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1797 = 10'h205 == io_inputs_1 ? 7'h0 : _GEN_1796; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1798 = 10'h206 == io_inputs_1 ? 7'h0 : _GEN_1797; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1799 = 10'h207 == io_inputs_1 ? 7'h0 : _GEN_1798; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1800 = 10'h208 == io_inputs_1 ? 7'h0 : _GEN_1799; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1801 = 10'h209 == io_inputs_1 ? 7'h0 : _GEN_1800; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1802 = 10'h20a == io_inputs_1 ? 7'h0 : _GEN_1801; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1803 = 10'h20b == io_inputs_1 ? 7'h0 : _GEN_1802; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1804 = 10'h20c == io_inputs_1 ? 7'h0 : _GEN_1803; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1805 = 10'h20d == io_inputs_1 ? 7'h0 : _GEN_1804; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1806 = 10'h20e == io_inputs_1 ? 7'h0 : _GEN_1805; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1807 = 10'h20f == io_inputs_1 ? 7'h0 : _GEN_1806; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1808 = 10'h210 == io_inputs_1 ? 7'h0 : _GEN_1807; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1809 = 10'h211 == io_inputs_1 ? 7'h0 : _GEN_1808; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1810 = 10'h212 == io_inputs_1 ? 7'h0 : _GEN_1809; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1811 = 10'h213 == io_inputs_1 ? 7'h0 : _GEN_1810; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1812 = 10'h214 == io_inputs_1 ? 7'h0 : _GEN_1811; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1813 = 10'h215 == io_inputs_1 ? 7'h0 : _GEN_1812; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1814 = 10'h216 == io_inputs_1 ? 7'h0 : _GEN_1813; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1815 = 10'h217 == io_inputs_1 ? 7'h0 : _GEN_1814; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1816 = 10'h218 == io_inputs_1 ? 7'h0 : _GEN_1815; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1817 = 10'h219 == io_inputs_1 ? 7'h0 : _GEN_1816; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1818 = 10'h21a == io_inputs_1 ? 7'h0 : _GEN_1817; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1819 = 10'h21b == io_inputs_1 ? 7'h0 : _GEN_1818; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1820 = 10'h21c == io_inputs_1 ? 7'h0 : _GEN_1819; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1821 = 10'h21d == io_inputs_1 ? 7'h0 : _GEN_1820; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1822 = 10'h21e == io_inputs_1 ? 7'h0 : _GEN_1821; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1823 = 10'h21f == io_inputs_1 ? 7'h0 : _GEN_1822; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1824 = 10'h220 == io_inputs_1 ? 7'h0 : _GEN_1823; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1825 = 10'h221 == io_inputs_1 ? 7'h0 : _GEN_1824; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1826 = 10'h222 == io_inputs_1 ? 7'h0 : _GEN_1825; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1827 = 10'h223 == io_inputs_1 ? 7'h0 : _GEN_1826; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1828 = 10'h224 == io_inputs_1 ? 7'h0 : _GEN_1827; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1829 = 10'h225 == io_inputs_1 ? 7'h0 : _GEN_1828; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1830 = 10'h226 == io_inputs_1 ? 7'h0 : _GEN_1829; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1831 = 10'h227 == io_inputs_1 ? 7'h0 : _GEN_1830; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1832 = 10'h228 == io_inputs_1 ? 7'h0 : _GEN_1831; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1833 = 10'h229 == io_inputs_1 ? 7'h0 : _GEN_1832; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1834 = 10'h22a == io_inputs_1 ? 7'h0 : _GEN_1833; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1835 = 10'h22b == io_inputs_1 ? 7'h0 : _GEN_1834; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1836 = 10'h22c == io_inputs_1 ? 7'h0 : _GEN_1835; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1837 = 10'h22d == io_inputs_1 ? 7'h0 : _GEN_1836; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1838 = 10'h22e == io_inputs_1 ? 7'h0 : _GEN_1837; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1839 = 10'h22f == io_inputs_1 ? 7'h0 : _GEN_1838; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1840 = 10'h230 == io_inputs_1 ? 7'h0 : _GEN_1839; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1841 = 10'h231 == io_inputs_1 ? 7'h0 : _GEN_1840; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1842 = 10'h232 == io_inputs_1 ? 7'h0 : _GEN_1841; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1843 = 10'h233 == io_inputs_1 ? 7'h0 : _GEN_1842; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1844 = 10'h234 == io_inputs_1 ? 7'h0 : _GEN_1843; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1845 = 10'h235 == io_inputs_1 ? 7'h0 : _GEN_1844; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1846 = 10'h236 == io_inputs_1 ? 7'h0 : _GEN_1845; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1847 = 10'h237 == io_inputs_1 ? 7'h0 : _GEN_1846; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1848 = 10'h238 == io_inputs_1 ? 7'h0 : _GEN_1847; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1849 = 10'h239 == io_inputs_1 ? 7'h0 : _GEN_1848; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1850 = 10'h23a == io_inputs_1 ? 7'h0 : _GEN_1849; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1851 = 10'h23b == io_inputs_1 ? 7'h0 : _GEN_1850; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1852 = 10'h23c == io_inputs_1 ? 7'h0 : _GEN_1851; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1853 = 10'h23d == io_inputs_1 ? 7'h0 : _GEN_1852; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1854 = 10'h23e == io_inputs_1 ? 7'h0 : _GEN_1853; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1855 = 10'h23f == io_inputs_1 ? 7'h0 : _GEN_1854; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1856 = 10'h240 == io_inputs_1 ? 7'h0 : _GEN_1855; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1857 = 10'h241 == io_inputs_1 ? 7'h0 : _GEN_1856; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1858 = 10'h242 == io_inputs_1 ? 7'h0 : _GEN_1857; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1859 = 10'h243 == io_inputs_1 ? 7'h0 : _GEN_1858; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1860 = 10'h244 == io_inputs_1 ? 7'h0 : _GEN_1859; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1861 = 10'h245 == io_inputs_1 ? 7'h0 : _GEN_1860; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1862 = 10'h246 == io_inputs_1 ? 7'h0 : _GEN_1861; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1863 = 10'h247 == io_inputs_1 ? 7'h0 : _GEN_1862; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1864 = 10'h248 == io_inputs_1 ? 7'h0 : _GEN_1863; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1865 = 10'h249 == io_inputs_1 ? 7'h0 : _GEN_1864; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1866 = 10'h24a == io_inputs_1 ? 7'h0 : _GEN_1865; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1867 = 10'h24b == io_inputs_1 ? 7'h0 : _GEN_1866; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1868 = 10'h24c == io_inputs_1 ? 7'h0 : _GEN_1867; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1869 = 10'h24d == io_inputs_1 ? 7'h0 : _GEN_1868; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1870 = 10'h24e == io_inputs_1 ? 7'h0 : _GEN_1869; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1871 = 10'h24f == io_inputs_1 ? 7'h0 : _GEN_1870; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1872 = 10'h250 == io_inputs_1 ? 7'h0 : _GEN_1871; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1873 = 10'h251 == io_inputs_1 ? 7'h0 : _GEN_1872; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1874 = 10'h252 == io_inputs_1 ? 7'h0 : _GEN_1873; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1875 = 10'h253 == io_inputs_1 ? 7'h0 : _GEN_1874; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1876 = 10'h254 == io_inputs_1 ? 7'h0 : _GEN_1875; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1877 = 10'h255 == io_inputs_1 ? 7'h0 : _GEN_1876; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1878 = 10'h256 == io_inputs_1 ? 7'h0 : _GEN_1877; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1879 = 10'h257 == io_inputs_1 ? 7'h0 : _GEN_1878; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1880 = 10'h258 == io_inputs_1 ? 7'h0 : _GEN_1879; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1881 = 10'h259 == io_inputs_1 ? 7'h0 : _GEN_1880; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1882 = 10'h25a == io_inputs_1 ? 7'h0 : _GEN_1881; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1883 = 10'h25b == io_inputs_1 ? 7'h0 : _GEN_1882; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1884 = 10'h25c == io_inputs_1 ? 7'h0 : _GEN_1883; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1885 = 10'h25d == io_inputs_1 ? 7'h0 : _GEN_1884; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1886 = 10'h25e == io_inputs_1 ? 7'h0 : _GEN_1885; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1887 = 10'h25f == io_inputs_1 ? 7'h0 : _GEN_1886; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1888 = 10'h260 == io_inputs_1 ? 7'h0 : _GEN_1887; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1889 = 10'h261 == io_inputs_1 ? 7'h0 : _GEN_1888; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1890 = 10'h262 == io_inputs_1 ? 7'h0 : _GEN_1889; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1891 = 10'h263 == io_inputs_1 ? 7'h0 : _GEN_1890; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1892 = 10'h264 == io_inputs_1 ? 7'h0 : _GEN_1891; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1893 = 10'h265 == io_inputs_1 ? 7'h0 : _GEN_1892; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1894 = 10'h266 == io_inputs_1 ? 7'h0 : _GEN_1893; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1895 = 10'h267 == io_inputs_1 ? 7'h0 : _GEN_1894; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1896 = 10'h268 == io_inputs_1 ? 7'h0 : _GEN_1895; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1897 = 10'h269 == io_inputs_1 ? 7'h0 : _GEN_1896; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1898 = 10'h26a == io_inputs_1 ? 7'h0 : _GEN_1897; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1899 = 10'h26b == io_inputs_1 ? 7'h0 : _GEN_1898; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1900 = 10'h26c == io_inputs_1 ? 7'h0 : _GEN_1899; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1901 = 10'h26d == io_inputs_1 ? 7'h0 : _GEN_1900; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1902 = 10'h26e == io_inputs_1 ? 7'h0 : _GEN_1901; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1903 = 10'h26f == io_inputs_1 ? 7'h0 : _GEN_1902; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1904 = 10'h270 == io_inputs_1 ? 7'h0 : _GEN_1903; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1905 = 10'h271 == io_inputs_1 ? 7'h0 : _GEN_1904; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1906 = 10'h272 == io_inputs_1 ? 7'h0 : _GEN_1905; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1907 = 10'h273 == io_inputs_1 ? 7'h0 : _GEN_1906; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1908 = 10'h274 == io_inputs_1 ? 7'h0 : _GEN_1907; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1909 = 10'h275 == io_inputs_1 ? 7'h0 : _GEN_1908; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1910 = 10'h276 == io_inputs_1 ? 7'h0 : _GEN_1909; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1911 = 10'h277 == io_inputs_1 ? 7'h0 : _GEN_1910; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1912 = 10'h278 == io_inputs_1 ? 7'h0 : _GEN_1911; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1913 = 10'h279 == io_inputs_1 ? 7'h0 : _GEN_1912; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1914 = 10'h27a == io_inputs_1 ? 7'h0 : _GEN_1913; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1915 = 10'h27b == io_inputs_1 ? 7'h0 : _GEN_1914; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1916 = 10'h27c == io_inputs_1 ? 7'h0 : _GEN_1915; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1917 = 10'h27d == io_inputs_1 ? 7'h0 : _GEN_1916; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1918 = 10'h27e == io_inputs_1 ? 7'h0 : _GEN_1917; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1919 = 10'h27f == io_inputs_1 ? 7'h0 : _GEN_1918; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1920 = 10'h280 == io_inputs_1 ? 7'h0 : _GEN_1919; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1921 = 10'h281 == io_inputs_1 ? 7'h0 : _GEN_1920; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1922 = 10'h282 == io_inputs_1 ? 7'h0 : _GEN_1921; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1923 = 10'h283 == io_inputs_1 ? 7'h0 : _GEN_1922; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1924 = 10'h284 == io_inputs_1 ? 7'h0 : _GEN_1923; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1925 = 10'h285 == io_inputs_1 ? 7'h0 : _GEN_1924; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1926 = 10'h286 == io_inputs_1 ? 7'h0 : _GEN_1925; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1927 = 10'h287 == io_inputs_1 ? 7'h0 : _GEN_1926; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1928 = 10'h288 == io_inputs_1 ? 7'h0 : _GEN_1927; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1929 = 10'h289 == io_inputs_1 ? 7'h0 : _GEN_1928; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1930 = 10'h28a == io_inputs_1 ? 7'h0 : _GEN_1929; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1931 = 10'h28b == io_inputs_1 ? 7'h0 : _GEN_1930; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1932 = 10'h28c == io_inputs_1 ? 7'h0 : _GEN_1931; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1933 = 10'h28d == io_inputs_1 ? 7'h0 : _GEN_1932; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1934 = 10'h28e == io_inputs_1 ? 7'h0 : _GEN_1933; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1935 = 10'h28f == io_inputs_1 ? 7'h0 : _GEN_1934; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1936 = 10'h290 == io_inputs_1 ? 7'h0 : _GEN_1935; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1937 = 10'h291 == io_inputs_1 ? 7'h0 : _GEN_1936; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1938 = 10'h292 == io_inputs_1 ? 7'h0 : _GEN_1937; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1939 = 10'h293 == io_inputs_1 ? 7'h0 : _GEN_1938; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1940 = 10'h294 == io_inputs_1 ? 7'h0 : _GEN_1939; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1941 = 10'h295 == io_inputs_1 ? 7'h0 : _GEN_1940; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1942 = 10'h296 == io_inputs_1 ? 7'h0 : _GEN_1941; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1943 = 10'h297 == io_inputs_1 ? 7'h0 : _GEN_1942; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1944 = 10'h298 == io_inputs_1 ? 7'h0 : _GEN_1943; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1945 = 10'h299 == io_inputs_1 ? 7'h0 : _GEN_1944; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1946 = 10'h29a == io_inputs_1 ? 7'h0 : _GEN_1945; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1947 = 10'h29b == io_inputs_1 ? 7'h0 : _GEN_1946; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1948 = 10'h29c == io_inputs_1 ? 7'h0 : _GEN_1947; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1949 = 10'h29d == io_inputs_1 ? 7'h0 : _GEN_1948; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1950 = 10'h29e == io_inputs_1 ? 7'h0 : _GEN_1949; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1951 = 10'h29f == io_inputs_1 ? 7'h0 : _GEN_1950; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1952 = 10'h2a0 == io_inputs_1 ? 7'h0 : _GEN_1951; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1953 = 10'h2a1 == io_inputs_1 ? 7'h0 : _GEN_1952; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1954 = 10'h2a2 == io_inputs_1 ? 7'h0 : _GEN_1953; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1955 = 10'h2a3 == io_inputs_1 ? 7'h0 : _GEN_1954; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1956 = 10'h2a4 == io_inputs_1 ? 7'h0 : _GEN_1955; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1957 = 10'h2a5 == io_inputs_1 ? 7'h0 : _GEN_1956; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1958 = 10'h2a6 == io_inputs_1 ? 7'h0 : _GEN_1957; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1959 = 10'h2a7 == io_inputs_1 ? 7'h0 : _GEN_1958; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1960 = 10'h2a8 == io_inputs_1 ? 7'h0 : _GEN_1959; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1961 = 10'h2a9 == io_inputs_1 ? 7'h0 : _GEN_1960; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1962 = 10'h2aa == io_inputs_1 ? 7'h0 : _GEN_1961; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1963 = 10'h2ab == io_inputs_1 ? 7'h0 : _GEN_1962; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1964 = 10'h2ac == io_inputs_1 ? 7'h0 : _GEN_1963; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1965 = 10'h2ad == io_inputs_1 ? 7'h0 : _GEN_1964; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1966 = 10'h2ae == io_inputs_1 ? 7'h0 : _GEN_1965; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1967 = 10'h2af == io_inputs_1 ? 7'h0 : _GEN_1966; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1968 = 10'h2b0 == io_inputs_1 ? 7'h0 : _GEN_1967; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1969 = 10'h2b1 == io_inputs_1 ? 7'h0 : _GEN_1968; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1970 = 10'h2b2 == io_inputs_1 ? 7'h0 : _GEN_1969; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1971 = 10'h2b3 == io_inputs_1 ? 7'h0 : _GEN_1970; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1972 = 10'h2b4 == io_inputs_1 ? 7'h0 : _GEN_1971; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1973 = 10'h2b5 == io_inputs_1 ? 7'h0 : _GEN_1972; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1974 = 10'h2b6 == io_inputs_1 ? 7'h0 : _GEN_1973; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1975 = 10'h2b7 == io_inputs_1 ? 7'h0 : _GEN_1974; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1976 = 10'h2b8 == io_inputs_1 ? 7'h0 : _GEN_1975; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1977 = 10'h2b9 == io_inputs_1 ? 7'h0 : _GEN_1976; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1978 = 10'h2ba == io_inputs_1 ? 7'h0 : _GEN_1977; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1979 = 10'h2bb == io_inputs_1 ? 7'h0 : _GEN_1978; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1980 = 10'h2bc == io_inputs_1 ? 7'h0 : _GEN_1979; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1981 = 10'h2bd == io_inputs_1 ? 7'h0 : _GEN_1980; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1982 = 10'h2be == io_inputs_1 ? 7'h0 : _GEN_1981; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1983 = 10'h2bf == io_inputs_1 ? 7'h0 : _GEN_1982; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1984 = 10'h2c0 == io_inputs_1 ? 7'h0 : _GEN_1983; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1985 = 10'h2c1 == io_inputs_1 ? 7'h0 : _GEN_1984; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1986 = 10'h2c2 == io_inputs_1 ? 7'h0 : _GEN_1985; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1987 = 10'h2c3 == io_inputs_1 ? 7'h0 : _GEN_1986; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1988 = 10'h2c4 == io_inputs_1 ? 7'h0 : _GEN_1987; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1989 = 10'h2c5 == io_inputs_1 ? 7'h0 : _GEN_1988; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1990 = 10'h2c6 == io_inputs_1 ? 7'h0 : _GEN_1989; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1991 = 10'h2c7 == io_inputs_1 ? 7'h0 : _GEN_1990; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1992 = 10'h2c8 == io_inputs_1 ? 7'h0 : _GEN_1991; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1993 = 10'h2c9 == io_inputs_1 ? 7'h0 : _GEN_1992; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1994 = 10'h2ca == io_inputs_1 ? 7'h0 : _GEN_1993; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1995 = 10'h2cb == io_inputs_1 ? 7'h0 : _GEN_1994; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1996 = 10'h2cc == io_inputs_1 ? 7'h0 : _GEN_1995; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1997 = 10'h2cd == io_inputs_1 ? 7'h0 : _GEN_1996; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1998 = 10'h2ce == io_inputs_1 ? 7'h0 : _GEN_1997; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_1999 = 10'h2cf == io_inputs_1 ? 7'h0 : _GEN_1998; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2000 = 10'h2d0 == io_inputs_1 ? 7'h0 : _GEN_1999; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2001 = 10'h2d1 == io_inputs_1 ? 7'h0 : _GEN_2000; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2002 = 10'h2d2 == io_inputs_1 ? 7'h0 : _GEN_2001; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2003 = 10'h2d3 == io_inputs_1 ? 7'h0 : _GEN_2002; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2004 = 10'h2d4 == io_inputs_1 ? 7'h0 : _GEN_2003; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2005 = 10'h2d5 == io_inputs_1 ? 7'h0 : _GEN_2004; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2006 = 10'h2d6 == io_inputs_1 ? 7'h0 : _GEN_2005; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2007 = 10'h2d7 == io_inputs_1 ? 7'h0 : _GEN_2006; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2008 = 10'h2d8 == io_inputs_1 ? 7'h0 : _GEN_2007; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2009 = 10'h2d9 == io_inputs_1 ? 7'h0 : _GEN_2008; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2010 = 10'h2da == io_inputs_1 ? 7'h0 : _GEN_2009; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2011 = 10'h2db == io_inputs_1 ? 7'h0 : _GEN_2010; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2012 = 10'h2dc == io_inputs_1 ? 7'h0 : _GEN_2011; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2013 = 10'h2dd == io_inputs_1 ? 7'h0 : _GEN_2012; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2014 = 10'h2de == io_inputs_1 ? 7'h0 : _GEN_2013; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2015 = 10'h2df == io_inputs_1 ? 7'h0 : _GEN_2014; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2016 = 10'h2e0 == io_inputs_1 ? 7'h0 : _GEN_2015; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2017 = 10'h2e1 == io_inputs_1 ? 7'h0 : _GEN_2016; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2018 = 10'h2e2 == io_inputs_1 ? 7'h0 : _GEN_2017; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2019 = 10'h2e3 == io_inputs_1 ? 7'h0 : _GEN_2018; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2020 = 10'h2e4 == io_inputs_1 ? 7'h0 : _GEN_2019; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2021 = 10'h2e5 == io_inputs_1 ? 7'h0 : _GEN_2020; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2022 = 10'h2e6 == io_inputs_1 ? 7'h0 : _GEN_2021; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2023 = 10'h2e7 == io_inputs_1 ? 7'h0 : _GEN_2022; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2024 = 10'h2e8 == io_inputs_1 ? 7'h0 : _GEN_2023; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2025 = 10'h2e9 == io_inputs_1 ? 7'h0 : _GEN_2024; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2026 = 10'h2ea == io_inputs_1 ? 7'h0 : _GEN_2025; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2027 = 10'h2eb == io_inputs_1 ? 7'h0 : _GEN_2026; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2028 = 10'h2ec == io_inputs_1 ? 7'h0 : _GEN_2027; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2029 = 10'h2ed == io_inputs_1 ? 7'h0 : _GEN_2028; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2030 = 10'h2ee == io_inputs_1 ? 7'h0 : _GEN_2029; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2031 = 10'h2ef == io_inputs_1 ? 7'h0 : _GEN_2030; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2032 = 10'h2f0 == io_inputs_1 ? 7'h0 : _GEN_2031; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2033 = 10'h2f1 == io_inputs_1 ? 7'h0 : _GEN_2032; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2034 = 10'h2f2 == io_inputs_1 ? 7'h0 : _GEN_2033; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2035 = 10'h2f3 == io_inputs_1 ? 7'h0 : _GEN_2034; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2036 = 10'h2f4 == io_inputs_1 ? 7'h0 : _GEN_2035; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2037 = 10'h2f5 == io_inputs_1 ? 7'h0 : _GEN_2036; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2038 = 10'h2f6 == io_inputs_1 ? 7'h0 : _GEN_2037; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2039 = 10'h2f7 == io_inputs_1 ? 7'h0 : _GEN_2038; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2040 = 10'h2f8 == io_inputs_1 ? 7'h0 : _GEN_2039; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2041 = 10'h2f9 == io_inputs_1 ? 7'h0 : _GEN_2040; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2042 = 10'h2fa == io_inputs_1 ? 7'h0 : _GEN_2041; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2043 = 10'h2fb == io_inputs_1 ? 7'h0 : _GEN_2042; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2044 = 10'h2fc == io_inputs_1 ? 7'h0 : _GEN_2043; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2045 = 10'h2fd == io_inputs_1 ? 7'h0 : _GEN_2044; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2046 = 10'h2fe == io_inputs_1 ? 7'h0 : _GEN_2045; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2047 = 10'h2ff == io_inputs_1 ? 7'h0 : _GEN_2046; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2048 = 10'h300 == io_inputs_1 ? 7'h0 : _GEN_2047; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2049 = 10'h301 == io_inputs_1 ? 7'h0 : _GEN_2048; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2050 = 10'h302 == io_inputs_1 ? 7'h0 : _GEN_2049; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2051 = 10'h303 == io_inputs_1 ? 7'h0 : _GEN_2050; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2052 = 10'h304 == io_inputs_1 ? 7'h0 : _GEN_2051; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2053 = 10'h305 == io_inputs_1 ? 7'h0 : _GEN_2052; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2054 = 10'h306 == io_inputs_1 ? 7'h0 : _GEN_2053; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2055 = 10'h307 == io_inputs_1 ? 7'h0 : _GEN_2054; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2056 = 10'h308 == io_inputs_1 ? 7'h0 : _GEN_2055; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2057 = 10'h309 == io_inputs_1 ? 7'h0 : _GEN_2056; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2058 = 10'h30a == io_inputs_1 ? 7'h0 : _GEN_2057; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2059 = 10'h30b == io_inputs_1 ? 7'h0 : _GEN_2058; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2060 = 10'h30c == io_inputs_1 ? 7'h0 : _GEN_2059; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2061 = 10'h30d == io_inputs_1 ? 7'h0 : _GEN_2060; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2062 = 10'h30e == io_inputs_1 ? 7'h0 : _GEN_2061; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2063 = 10'h30f == io_inputs_1 ? 7'h0 : _GEN_2062; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2064 = 10'h310 == io_inputs_1 ? 7'h0 : _GEN_2063; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2065 = 10'h311 == io_inputs_1 ? 7'h0 : _GEN_2064; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2066 = 10'h312 == io_inputs_1 ? 7'h0 : _GEN_2065; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2067 = 10'h313 == io_inputs_1 ? 7'h0 : _GEN_2066; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2068 = 10'h314 == io_inputs_1 ? 7'h0 : _GEN_2067; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2069 = 10'h315 == io_inputs_1 ? 7'h0 : _GEN_2068; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2070 = 10'h316 == io_inputs_1 ? 7'h0 : _GEN_2069; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2071 = 10'h317 == io_inputs_1 ? 7'h0 : _GEN_2070; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2072 = 10'h318 == io_inputs_1 ? 7'h0 : _GEN_2071; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2073 = 10'h319 == io_inputs_1 ? 7'h0 : _GEN_2072; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2074 = 10'h31a == io_inputs_1 ? 7'h0 : _GEN_2073; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2075 = 10'h31b == io_inputs_1 ? 7'h0 : _GEN_2074; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2076 = 10'h31c == io_inputs_1 ? 7'h0 : _GEN_2075; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2077 = 10'h31d == io_inputs_1 ? 7'h0 : _GEN_2076; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2078 = 10'h31e == io_inputs_1 ? 7'h0 : _GEN_2077; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2079 = 10'h31f == io_inputs_1 ? 7'h0 : _GEN_2078; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2080 = 10'h320 == io_inputs_1 ? 7'h0 : _GEN_2079; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2081 = 10'h321 == io_inputs_1 ? 7'h0 : _GEN_2080; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2082 = 10'h322 == io_inputs_1 ? 7'h0 : _GEN_2081; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2083 = 10'h323 == io_inputs_1 ? 7'h0 : _GEN_2082; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2084 = 10'h324 == io_inputs_1 ? 7'h0 : _GEN_2083; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2085 = 10'h325 == io_inputs_1 ? 7'h0 : _GEN_2084; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2086 = 10'h326 == io_inputs_1 ? 7'h0 : _GEN_2085; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2087 = 10'h327 == io_inputs_1 ? 7'h0 : _GEN_2086; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2088 = 10'h328 == io_inputs_1 ? 7'h0 : _GEN_2087; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2089 = 10'h329 == io_inputs_1 ? 7'h0 : _GEN_2088; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2090 = 10'h32a == io_inputs_1 ? 7'h0 : _GEN_2089; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2091 = 10'h32b == io_inputs_1 ? 7'h0 : _GEN_2090; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2092 = 10'h32c == io_inputs_1 ? 7'h0 : _GEN_2091; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2093 = 10'h32d == io_inputs_1 ? 7'h0 : _GEN_2092; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2094 = 10'h32e == io_inputs_1 ? 7'h0 : _GEN_2093; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2095 = 10'h32f == io_inputs_1 ? 7'h0 : _GEN_2094; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2096 = 10'h330 == io_inputs_1 ? 7'h0 : _GEN_2095; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2097 = 10'h331 == io_inputs_1 ? 7'h0 : _GEN_2096; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2098 = 10'h332 == io_inputs_1 ? 7'h0 : _GEN_2097; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2099 = 10'h333 == io_inputs_1 ? 7'h0 : _GEN_2098; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2100 = 10'h334 == io_inputs_1 ? 7'h0 : _GEN_2099; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2101 = 10'h335 == io_inputs_1 ? 7'h0 : _GEN_2100; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2102 = 10'h336 == io_inputs_1 ? 7'h0 : _GEN_2101; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2103 = 10'h337 == io_inputs_1 ? 7'h0 : _GEN_2102; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2104 = 10'h338 == io_inputs_1 ? 7'h0 : _GEN_2103; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2105 = 10'h339 == io_inputs_1 ? 7'h0 : _GEN_2104; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2106 = 10'h33a == io_inputs_1 ? 7'h0 : _GEN_2105; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2107 = 10'h33b == io_inputs_1 ? 7'h0 : _GEN_2106; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2108 = 10'h33c == io_inputs_1 ? 7'h0 : _GEN_2107; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2109 = 10'h33d == io_inputs_1 ? 7'h0 : _GEN_2108; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2110 = 10'h33e == io_inputs_1 ? 7'h0 : _GEN_2109; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2111 = 10'h33f == io_inputs_1 ? 7'h0 : _GEN_2110; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2112 = 10'h340 == io_inputs_1 ? 7'h0 : _GEN_2111; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2113 = 10'h341 == io_inputs_1 ? 7'h0 : _GEN_2112; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2114 = 10'h342 == io_inputs_1 ? 7'h0 : _GEN_2113; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2115 = 10'h343 == io_inputs_1 ? 7'h0 : _GEN_2114; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2116 = 10'h344 == io_inputs_1 ? 7'h0 : _GEN_2115; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2117 = 10'h345 == io_inputs_1 ? 7'h0 : _GEN_2116; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2118 = 10'h346 == io_inputs_1 ? 7'h0 : _GEN_2117; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2119 = 10'h347 == io_inputs_1 ? 7'h0 : _GEN_2118; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2120 = 10'h348 == io_inputs_1 ? 7'h0 : _GEN_2119; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2121 = 10'h349 == io_inputs_1 ? 7'h0 : _GEN_2120; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2122 = 10'h34a == io_inputs_1 ? 7'h0 : _GEN_2121; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2123 = 10'h34b == io_inputs_1 ? 7'h0 : _GEN_2122; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2124 = 10'h34c == io_inputs_1 ? 7'h0 : _GEN_2123; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2125 = 10'h34d == io_inputs_1 ? 7'h0 : _GEN_2124; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2126 = 10'h34e == io_inputs_1 ? 7'h0 : _GEN_2125; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2127 = 10'h34f == io_inputs_1 ? 7'h0 : _GEN_2126; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2128 = 10'h350 == io_inputs_1 ? 7'h0 : _GEN_2127; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2129 = 10'h351 == io_inputs_1 ? 7'h0 : _GEN_2128; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2130 = 10'h352 == io_inputs_1 ? 7'h0 : _GEN_2129; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2131 = 10'h353 == io_inputs_1 ? 7'h0 : _GEN_2130; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2132 = 10'h354 == io_inputs_1 ? 7'h0 : _GEN_2131; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2133 = 10'h355 == io_inputs_1 ? 7'h0 : _GEN_2132; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2134 = 10'h356 == io_inputs_1 ? 7'h0 : _GEN_2133; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2135 = 10'h357 == io_inputs_1 ? 7'h0 : _GEN_2134; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2136 = 10'h358 == io_inputs_1 ? 7'h0 : _GEN_2135; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2137 = 10'h359 == io_inputs_1 ? 7'h0 : _GEN_2136; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2138 = 10'h35a == io_inputs_1 ? 7'h0 : _GEN_2137; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2139 = 10'h35b == io_inputs_1 ? 7'h0 : _GEN_2138; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2140 = 10'h35c == io_inputs_1 ? 7'h0 : _GEN_2139; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2141 = 10'h35d == io_inputs_1 ? 7'h0 : _GEN_2140; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2142 = 10'h35e == io_inputs_1 ? 7'h0 : _GEN_2141; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2143 = 10'h35f == io_inputs_1 ? 7'h0 : _GEN_2142; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2144 = 10'h360 == io_inputs_1 ? 7'h0 : _GEN_2143; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2145 = 10'h361 == io_inputs_1 ? 7'h0 : _GEN_2144; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2146 = 10'h362 == io_inputs_1 ? 7'h0 : _GEN_2145; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2147 = 10'h363 == io_inputs_1 ? 7'h0 : _GEN_2146; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2148 = 10'h364 == io_inputs_1 ? 7'h0 : _GEN_2147; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2149 = 10'h365 == io_inputs_1 ? 7'h0 : _GEN_2148; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2150 = 10'h366 == io_inputs_1 ? 7'h0 : _GEN_2149; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2151 = 10'h367 == io_inputs_1 ? 7'h0 : _GEN_2150; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2152 = 10'h368 == io_inputs_1 ? 7'h0 : _GEN_2151; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2153 = 10'h369 == io_inputs_1 ? 7'h0 : _GEN_2152; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2154 = 10'h36a == io_inputs_1 ? 7'h0 : _GEN_2153; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2155 = 10'h36b == io_inputs_1 ? 7'h0 : _GEN_2154; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2156 = 10'h36c == io_inputs_1 ? 7'h0 : _GEN_2155; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2157 = 10'h36d == io_inputs_1 ? 7'h0 : _GEN_2156; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2158 = 10'h36e == io_inputs_1 ? 7'h0 : _GEN_2157; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2159 = 10'h36f == io_inputs_1 ? 7'h0 : _GEN_2158; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2160 = 10'h370 == io_inputs_1 ? 7'h0 : _GEN_2159; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2161 = 10'h371 == io_inputs_1 ? 7'h0 : _GEN_2160; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2162 = 10'h372 == io_inputs_1 ? 7'h0 : _GEN_2161; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2163 = 10'h373 == io_inputs_1 ? 7'h0 : _GEN_2162; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2164 = 10'h374 == io_inputs_1 ? 7'h0 : _GEN_2163; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2165 = 10'h375 == io_inputs_1 ? 7'h0 : _GEN_2164; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2166 = 10'h376 == io_inputs_1 ? 7'h0 : _GEN_2165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2167 = 10'h377 == io_inputs_1 ? 7'h0 : _GEN_2166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2168 = 10'h378 == io_inputs_1 ? 7'h0 : _GEN_2167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2169 = 10'h379 == io_inputs_1 ? 7'h0 : _GEN_2168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2170 = 10'h37a == io_inputs_1 ? 7'h0 : _GEN_2169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2171 = 10'h37b == io_inputs_1 ? 7'h0 : _GEN_2170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2172 = 10'h37c == io_inputs_1 ? 7'h0 : _GEN_2171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2173 = 10'h37d == io_inputs_1 ? 7'h0 : _GEN_2172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2174 = 10'h37e == io_inputs_1 ? 7'h0 : _GEN_2173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2175 = 10'h37f == io_inputs_1 ? 7'h0 : _GEN_2174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2176 = 10'h380 == io_inputs_1 ? 7'h0 : _GEN_2175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2177 = 10'h381 == io_inputs_1 ? 7'h0 : _GEN_2176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2178 = 10'h382 == io_inputs_1 ? 7'h0 : _GEN_2177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2179 = 10'h383 == io_inputs_1 ? 7'h0 : _GEN_2178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2180 = 10'h384 == io_inputs_1 ? 7'h0 : _GEN_2179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2181 = 10'h385 == io_inputs_1 ? 7'h0 : _GEN_2180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2182 = 10'h386 == io_inputs_1 ? 7'h0 : _GEN_2181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2183 = 10'h387 == io_inputs_1 ? 7'h0 : _GEN_2182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2184 = 10'h388 == io_inputs_1 ? 7'h0 : _GEN_2183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2185 = 10'h389 == io_inputs_1 ? 7'h0 : _GEN_2184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2186 = 10'h38a == io_inputs_1 ? 7'h0 : _GEN_2185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2187 = 10'h38b == io_inputs_1 ? 7'h0 : _GEN_2186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2188 = 10'h38c == io_inputs_1 ? 7'h0 : _GEN_2187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2189 = 10'h38d == io_inputs_1 ? 7'h0 : _GEN_2188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2190 = 10'h38e == io_inputs_1 ? 7'h0 : _GEN_2189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2191 = 10'h38f == io_inputs_1 ? 7'h0 : _GEN_2190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2192 = 10'h390 == io_inputs_1 ? 7'h0 : _GEN_2191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2193 = 10'h391 == io_inputs_1 ? 7'h0 : _GEN_2192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2194 = 10'h392 == io_inputs_1 ? 7'h0 : _GEN_2193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2195 = 10'h393 == io_inputs_1 ? 7'h0 : _GEN_2194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2196 = 10'h394 == io_inputs_1 ? 7'h0 : _GEN_2195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2197 = 10'h395 == io_inputs_1 ? 7'h0 : _GEN_2196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2198 = 10'h396 == io_inputs_1 ? 7'h0 : _GEN_2197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2199 = 10'h397 == io_inputs_1 ? 7'h0 : _GEN_2198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2200 = 10'h398 == io_inputs_1 ? 7'h0 : _GEN_2199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2201 = 10'h399 == io_inputs_1 ? 7'h0 : _GEN_2200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2202 = 10'h39a == io_inputs_1 ? 7'h0 : _GEN_2201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2203 = 10'h39b == io_inputs_1 ? 7'h0 : _GEN_2202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2204 = 10'h39c == io_inputs_1 ? 7'h0 : _GEN_2203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2205 = 10'h39d == io_inputs_1 ? 7'h0 : _GEN_2204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2206 = 10'h39e == io_inputs_1 ? 7'h0 : _GEN_2205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2207 = 10'h39f == io_inputs_1 ? 7'h0 : _GEN_2206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2208 = 10'h3a0 == io_inputs_1 ? 7'h0 : _GEN_2207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2209 = 10'h3a1 == io_inputs_1 ? 7'h0 : _GEN_2208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2210 = 10'h3a2 == io_inputs_1 ? 7'h0 : _GEN_2209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2211 = 10'h3a3 == io_inputs_1 ? 7'h0 : _GEN_2210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2212 = 10'h3a4 == io_inputs_1 ? 7'h0 : _GEN_2211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2213 = 10'h3a5 == io_inputs_1 ? 7'h0 : _GEN_2212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2214 = 10'h3a6 == io_inputs_1 ? 7'h0 : _GEN_2213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2215 = 10'h3a7 == io_inputs_1 ? 7'h0 : _GEN_2214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2216 = 10'h3a8 == io_inputs_1 ? 7'h0 : _GEN_2215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2217 = 10'h3a9 == io_inputs_1 ? 7'h0 : _GEN_2216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2218 = 10'h3aa == io_inputs_1 ? 7'h0 : _GEN_2217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2219 = 10'h3ab == io_inputs_1 ? 7'h0 : _GEN_2218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2220 = 10'h3ac == io_inputs_1 ? 7'h0 : _GEN_2219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2221 = 10'h3ad == io_inputs_1 ? 7'h0 : _GEN_2220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2222 = 10'h3ae == io_inputs_1 ? 7'h0 : _GEN_2221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2223 = 10'h3af == io_inputs_1 ? 7'h0 : _GEN_2222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2224 = 10'h3b0 == io_inputs_1 ? 7'h0 : _GEN_2223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2225 = 10'h3b1 == io_inputs_1 ? 7'h0 : _GEN_2224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2226 = 10'h3b2 == io_inputs_1 ? 7'h0 : _GEN_2225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2227 = 10'h3b3 == io_inputs_1 ? 7'h0 : _GEN_2226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2228 = 10'h3b4 == io_inputs_1 ? 7'h0 : _GEN_2227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2229 = 10'h3b5 == io_inputs_1 ? 7'h0 : _GEN_2228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2230 = 10'h3b6 == io_inputs_1 ? 7'h0 : _GEN_2229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2231 = 10'h3b7 == io_inputs_1 ? 7'h0 : _GEN_2230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2232 = 10'h3b8 == io_inputs_1 ? 7'h0 : _GEN_2231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2233 = 10'h3b9 == io_inputs_1 ? 7'h0 : _GEN_2232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2234 = 10'h3ba == io_inputs_1 ? 7'h0 : _GEN_2233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2235 = 10'h3bb == io_inputs_1 ? 7'h0 : _GEN_2234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2236 = 10'h3bc == io_inputs_1 ? 7'h0 : _GEN_2235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2237 = 10'h3bd == io_inputs_1 ? 7'h0 : _GEN_2236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2238 = 10'h3be == io_inputs_1 ? 7'h0 : _GEN_2237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2239 = 10'h3bf == io_inputs_1 ? 7'h0 : _GEN_2238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2240 = 10'h3c0 == io_inputs_1 ? 7'h0 : _GEN_2239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2241 = 10'h3c1 == io_inputs_1 ? 7'h0 : _GEN_2240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2242 = 10'h3c2 == io_inputs_1 ? 7'h0 : _GEN_2241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2243 = 10'h3c3 == io_inputs_1 ? 7'h0 : _GEN_2242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2244 = 10'h3c4 == io_inputs_1 ? 7'h0 : _GEN_2243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2245 = 10'h3c5 == io_inputs_1 ? 7'h0 : _GEN_2244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2246 = 10'h3c6 == io_inputs_1 ? 7'h0 : _GEN_2245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2247 = 10'h3c7 == io_inputs_1 ? 7'h0 : _GEN_2246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2248 = 10'h3c8 == io_inputs_1 ? 7'h0 : _GEN_2247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2249 = 10'h3c9 == io_inputs_1 ? 7'h0 : _GEN_2248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2250 = 10'h3ca == io_inputs_1 ? 7'h0 : _GEN_2249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2251 = 10'h3cb == io_inputs_1 ? 7'h0 : _GEN_2250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2252 = 10'h3cc == io_inputs_1 ? 7'h0 : _GEN_2251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2253 = 10'h3cd == io_inputs_1 ? 7'h0 : _GEN_2252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2254 = 10'h3ce == io_inputs_1 ? 7'h0 : _GEN_2253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2255 = 10'h3cf == io_inputs_1 ? 7'h0 : _GEN_2254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2256 = 10'h3d0 == io_inputs_1 ? 7'h0 : _GEN_2255; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2257 = 10'h3d1 == io_inputs_1 ? 7'h0 : _GEN_2256; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2258 = 10'h3d2 == io_inputs_1 ? 7'h0 : _GEN_2257; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2259 = 10'h3d3 == io_inputs_1 ? 7'h0 : _GEN_2258; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2260 = 10'h3d4 == io_inputs_1 ? 7'h0 : _GEN_2259; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2261 = 10'h3d5 == io_inputs_1 ? 7'h0 : _GEN_2260; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2262 = 10'h3d6 == io_inputs_1 ? 7'h0 : _GEN_2261; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2263 = 10'h3d7 == io_inputs_1 ? 7'h0 : _GEN_2262; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2264 = 10'h3d8 == io_inputs_1 ? 7'h0 : _GEN_2263; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2265 = 10'h3d9 == io_inputs_1 ? 7'h0 : _GEN_2264; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2266 = 10'h3da == io_inputs_1 ? 7'h0 : _GEN_2265; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2267 = 10'h3db == io_inputs_1 ? 7'h0 : _GEN_2266; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2268 = 10'h3dc == io_inputs_1 ? 7'h0 : _GEN_2267; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2269 = 10'h3dd == io_inputs_1 ? 7'h0 : _GEN_2268; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2270 = 10'h3de == io_inputs_1 ? 7'h0 : _GEN_2269; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2271 = 10'h3df == io_inputs_1 ? 7'h0 : _GEN_2270; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2272 = 10'h3e0 == io_inputs_1 ? 7'h0 : _GEN_2271; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2273 = 10'h3e1 == io_inputs_1 ? 7'h0 : _GEN_2272; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2274 = 10'h3e2 == io_inputs_1 ? 7'h0 : _GEN_2273; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2275 = 10'h3e3 == io_inputs_1 ? 7'h0 : _GEN_2274; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2276 = 10'h3e4 == io_inputs_1 ? 7'h0 : _GEN_2275; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2277 = 10'h3e5 == io_inputs_1 ? 7'h0 : _GEN_2276; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2278 = 10'h3e6 == io_inputs_1 ? 7'h0 : _GEN_2277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2279 = 10'h3e7 == io_inputs_1 ? 7'h0 : _GEN_2278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2280 = 10'h3e8 == io_inputs_1 ? 7'h0 : _GEN_2279; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2281 = 10'h3e9 == io_inputs_1 ? 7'h0 : _GEN_2280; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2282 = 10'h3ea == io_inputs_1 ? 7'h0 : _GEN_2281; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2283 = 10'h3eb == io_inputs_1 ? 7'h0 : _GEN_2282; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2284 = 10'h3ec == io_inputs_1 ? 7'h0 : _GEN_2283; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2285 = 10'h3ed == io_inputs_1 ? 7'h0 : _GEN_2284; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2286 = 10'h3ee == io_inputs_1 ? 7'h0 : _GEN_2285; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2287 = 10'h3ef == io_inputs_1 ? 7'h0 : _GEN_2286; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2288 = 10'h3f0 == io_inputs_1 ? 7'h0 : _GEN_2287; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2289 = 10'h3f1 == io_inputs_1 ? 7'h0 : _GEN_2288; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2290 = 10'h3f2 == io_inputs_1 ? 7'h0 : _GEN_2289; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2291 = 10'h3f3 == io_inputs_1 ? 7'h0 : _GEN_2290; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2292 = 10'h3f4 == io_inputs_1 ? 7'h0 : _GEN_2291; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2293 = 10'h3f5 == io_inputs_1 ? 7'h0 : _GEN_2292; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2294 = 10'h3f6 == io_inputs_1 ? 7'h0 : _GEN_2293; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2295 = 10'h3f7 == io_inputs_1 ? 7'h0 : _GEN_2294; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2296 = 10'h3f8 == io_inputs_1 ? 7'h0 : _GEN_2295; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2297 = 10'h3f9 == io_inputs_1 ? 7'h0 : _GEN_2296; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2298 = 10'h3fa == io_inputs_1 ? 7'h0 : _GEN_2297; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2299 = 10'h3fb == io_inputs_1 ? 7'h0 : _GEN_2298; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2300 = 10'h3fc == io_inputs_1 ? 7'h0 : _GEN_2299; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2301 = 10'h3fd == io_inputs_1 ? 7'h0 : _GEN_2300; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2302 = 10'h3fe == io_inputs_1 ? 7'h0 : _GEN_2301; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2303 = 10'h3ff == io_inputs_1 ? 7'h0 : _GEN_2302; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2355 = 10'h33 == io_inputs_1 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2356 = 10'h34 == io_inputs_1 ? 7'h2 : _GEN_2355; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2357 = 10'h35 == io_inputs_1 ? 7'h3 : _GEN_2356; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2358 = 10'h36 == io_inputs_1 ? 7'h4 : _GEN_2357; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2359 = 10'h37 == io_inputs_1 ? 7'h5 : _GEN_2358; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2360 = 10'h38 == io_inputs_1 ? 7'h6 : _GEN_2359; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2361 = 10'h39 == io_inputs_1 ? 7'h7 : _GEN_2360; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2362 = 10'h3a == io_inputs_1 ? 7'h8 : _GEN_2361; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2363 = 10'h3b == io_inputs_1 ? 7'h9 : _GEN_2362; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2364 = 10'h3c == io_inputs_1 ? 7'ha : _GEN_2363; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2365 = 10'h3d == io_inputs_1 ? 7'hb : _GEN_2364; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2366 = 10'h3e == io_inputs_1 ? 7'hc : _GEN_2365; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2367 = 10'h3f == io_inputs_1 ? 7'hd : _GEN_2366; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2368 = 10'h40 == io_inputs_1 ? 7'he : _GEN_2367; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2369 = 10'h41 == io_inputs_1 ? 7'hf : _GEN_2368; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2370 = 10'h42 == io_inputs_1 ? 7'h10 : _GEN_2369; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2371 = 10'h43 == io_inputs_1 ? 7'h11 : _GEN_2370; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2372 = 10'h44 == io_inputs_1 ? 7'h12 : _GEN_2371; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2373 = 10'h45 == io_inputs_1 ? 7'h13 : _GEN_2372; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2374 = 10'h46 == io_inputs_1 ? 7'h14 : _GEN_2373; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2375 = 10'h47 == io_inputs_1 ? 7'h15 : _GEN_2374; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2376 = 10'h48 == io_inputs_1 ? 7'h16 : _GEN_2375; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2377 = 10'h49 == io_inputs_1 ? 7'h17 : _GEN_2376; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2378 = 10'h4a == io_inputs_1 ? 7'h18 : _GEN_2377; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2379 = 10'h4b == io_inputs_1 ? 7'h19 : _GEN_2378; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2380 = 10'h4c == io_inputs_1 ? 7'h1a : _GEN_2379; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2381 = 10'h4d == io_inputs_1 ? 7'h1b : _GEN_2380; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2382 = 10'h4e == io_inputs_1 ? 7'h1c : _GEN_2381; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2383 = 10'h4f == io_inputs_1 ? 7'h1d : _GEN_2382; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2384 = 10'h50 == io_inputs_1 ? 7'h1e : _GEN_2383; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2385 = 10'h51 == io_inputs_1 ? 7'h1f : _GEN_2384; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2386 = 10'h52 == io_inputs_1 ? 7'h20 : _GEN_2385; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2387 = 10'h53 == io_inputs_1 ? 7'h21 : _GEN_2386; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2388 = 10'h54 == io_inputs_1 ? 7'h22 : _GEN_2387; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2389 = 10'h55 == io_inputs_1 ? 7'h23 : _GEN_2388; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2390 = 10'h56 == io_inputs_1 ? 7'h24 : _GEN_2389; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2391 = 10'h57 == io_inputs_1 ? 7'h25 : _GEN_2390; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2392 = 10'h58 == io_inputs_1 ? 7'h26 : _GEN_2391; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2393 = 10'h59 == io_inputs_1 ? 7'h27 : _GEN_2392; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2394 = 10'h5a == io_inputs_1 ? 7'h28 : _GEN_2393; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2395 = 10'h5b == io_inputs_1 ? 7'h29 : _GEN_2394; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2396 = 10'h5c == io_inputs_1 ? 7'h2a : _GEN_2395; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2397 = 10'h5d == io_inputs_1 ? 7'h2b : _GEN_2396; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2398 = 10'h5e == io_inputs_1 ? 7'h2c : _GEN_2397; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2399 = 10'h5f == io_inputs_1 ? 7'h2d : _GEN_2398; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2400 = 10'h60 == io_inputs_1 ? 7'h2e : _GEN_2399; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2401 = 10'h61 == io_inputs_1 ? 7'h2f : _GEN_2400; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2402 = 10'h62 == io_inputs_1 ? 7'h30 : _GEN_2401; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2403 = 10'h63 == io_inputs_1 ? 7'h31 : _GEN_2402; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2404 = 10'h64 == io_inputs_1 ? 7'h32 : _GEN_2403; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2405 = 10'h65 == io_inputs_1 ? 7'h33 : _GEN_2404; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2406 = 10'h66 == io_inputs_1 ? 7'h34 : _GEN_2405; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2407 = 10'h67 == io_inputs_1 ? 7'h35 : _GEN_2406; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2408 = 10'h68 == io_inputs_1 ? 7'h36 : _GEN_2407; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2409 = 10'h69 == io_inputs_1 ? 7'h37 : _GEN_2408; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2410 = 10'h6a == io_inputs_1 ? 7'h38 : _GEN_2409; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2411 = 10'h6b == io_inputs_1 ? 7'h39 : _GEN_2410; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2412 = 10'h6c == io_inputs_1 ? 7'h3a : _GEN_2411; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2413 = 10'h6d == io_inputs_1 ? 7'h3b : _GEN_2412; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2414 = 10'h6e == io_inputs_1 ? 7'h3c : _GEN_2413; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2415 = 10'h6f == io_inputs_1 ? 7'h3d : _GEN_2414; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2416 = 10'h70 == io_inputs_1 ? 7'h3e : _GEN_2415; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2417 = 10'h71 == io_inputs_1 ? 7'h3f : _GEN_2416; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2418 = 10'h72 == io_inputs_1 ? 7'h40 : _GEN_2417; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2419 = 10'h73 == io_inputs_1 ? 7'h41 : _GEN_2418; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2420 = 10'h74 == io_inputs_1 ? 7'h42 : _GEN_2419; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2421 = 10'h75 == io_inputs_1 ? 7'h43 : _GEN_2420; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2422 = 10'h76 == io_inputs_1 ? 7'h44 : _GEN_2421; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2423 = 10'h77 == io_inputs_1 ? 7'h45 : _GEN_2422; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2424 = 10'h78 == io_inputs_1 ? 7'h46 : _GEN_2423; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2425 = 10'h79 == io_inputs_1 ? 7'h47 : _GEN_2424; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2426 = 10'h7a == io_inputs_1 ? 7'h48 : _GEN_2425; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2427 = 10'h7b == io_inputs_1 ? 7'h49 : _GEN_2426; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2428 = 10'h7c == io_inputs_1 ? 7'h4a : _GEN_2427; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2429 = 10'h7d == io_inputs_1 ? 7'h4b : _GEN_2428; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2430 = 10'h7e == io_inputs_1 ? 7'h4c : _GEN_2429; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2431 = 10'h7f == io_inputs_1 ? 7'h4d : _GEN_2430; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2432 = 10'h80 == io_inputs_1 ? 7'h4e : _GEN_2431; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2433 = 10'h81 == io_inputs_1 ? 7'h4f : _GEN_2432; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2434 = 10'h82 == io_inputs_1 ? 7'h50 : _GEN_2433; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2435 = 10'h83 == io_inputs_1 ? 7'h51 : _GEN_2434; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2436 = 10'h84 == io_inputs_1 ? 7'h52 : _GEN_2435; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2437 = 10'h85 == io_inputs_1 ? 7'h53 : _GEN_2436; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2438 = 10'h86 == io_inputs_1 ? 7'h54 : _GEN_2437; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2439 = 10'h87 == io_inputs_1 ? 7'h55 : _GEN_2438; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2440 = 10'h88 == io_inputs_1 ? 7'h56 : _GEN_2439; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2441 = 10'h89 == io_inputs_1 ? 7'h57 : _GEN_2440; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2442 = 10'h8a == io_inputs_1 ? 7'h58 : _GEN_2441; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2443 = 10'h8b == io_inputs_1 ? 7'h59 : _GEN_2442; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2444 = 10'h8c == io_inputs_1 ? 7'h5a : _GEN_2443; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2445 = 10'h8d == io_inputs_1 ? 7'h5b : _GEN_2444; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2446 = 10'h8e == io_inputs_1 ? 7'h5c : _GEN_2445; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2447 = 10'h8f == io_inputs_1 ? 7'h5d : _GEN_2446; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2448 = 10'h90 == io_inputs_1 ? 7'h5e : _GEN_2447; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2449 = 10'h91 == io_inputs_1 ? 7'h5f : _GEN_2448; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2450 = 10'h92 == io_inputs_1 ? 7'h60 : _GEN_2449; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2451 = 10'h93 == io_inputs_1 ? 7'h61 : _GEN_2450; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2452 = 10'h94 == io_inputs_1 ? 7'h62 : _GEN_2451; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2453 = 10'h95 == io_inputs_1 ? 7'h63 : _GEN_2452; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2454 = 10'h96 == io_inputs_1 ? 7'h64 : _GEN_2453; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2455 = 10'h97 == io_inputs_1 ? 7'h64 : _GEN_2454; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2456 = 10'h98 == io_inputs_1 ? 7'h64 : _GEN_2455; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2457 = 10'h99 == io_inputs_1 ? 7'h64 : _GEN_2456; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2458 = 10'h9a == io_inputs_1 ? 7'h64 : _GEN_2457; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2459 = 10'h9b == io_inputs_1 ? 7'h64 : _GEN_2458; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2460 = 10'h9c == io_inputs_1 ? 7'h64 : _GEN_2459; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2461 = 10'h9d == io_inputs_1 ? 7'h64 : _GEN_2460; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2462 = 10'h9e == io_inputs_1 ? 7'h64 : _GEN_2461; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2463 = 10'h9f == io_inputs_1 ? 7'h64 : _GEN_2462; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2464 = 10'ha0 == io_inputs_1 ? 7'h64 : _GEN_2463; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2465 = 10'ha1 == io_inputs_1 ? 7'h64 : _GEN_2464; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2466 = 10'ha2 == io_inputs_1 ? 7'h64 : _GEN_2465; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2467 = 10'ha3 == io_inputs_1 ? 7'h64 : _GEN_2466; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2468 = 10'ha4 == io_inputs_1 ? 7'h64 : _GEN_2467; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2469 = 10'ha5 == io_inputs_1 ? 7'h64 : _GEN_2468; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2470 = 10'ha6 == io_inputs_1 ? 7'h64 : _GEN_2469; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2471 = 10'ha7 == io_inputs_1 ? 7'h64 : _GEN_2470; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2472 = 10'ha8 == io_inputs_1 ? 7'h64 : _GEN_2471; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2473 = 10'ha9 == io_inputs_1 ? 7'h64 : _GEN_2472; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2474 = 10'haa == io_inputs_1 ? 7'h64 : _GEN_2473; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2475 = 10'hab == io_inputs_1 ? 7'h64 : _GEN_2474; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2476 = 10'hac == io_inputs_1 ? 7'h64 : _GEN_2475; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2477 = 10'had == io_inputs_1 ? 7'h64 : _GEN_2476; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2478 = 10'hae == io_inputs_1 ? 7'h64 : _GEN_2477; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2479 = 10'haf == io_inputs_1 ? 7'h64 : _GEN_2478; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2480 = 10'hb0 == io_inputs_1 ? 7'h64 : _GEN_2479; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2481 = 10'hb1 == io_inputs_1 ? 7'h64 : _GEN_2480; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2482 = 10'hb2 == io_inputs_1 ? 7'h64 : _GEN_2481; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2483 = 10'hb3 == io_inputs_1 ? 7'h64 : _GEN_2482; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2484 = 10'hb4 == io_inputs_1 ? 7'h64 : _GEN_2483; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2485 = 10'hb5 == io_inputs_1 ? 7'h64 : _GEN_2484; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2486 = 10'hb6 == io_inputs_1 ? 7'h64 : _GEN_2485; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2487 = 10'hb7 == io_inputs_1 ? 7'h64 : _GEN_2486; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2488 = 10'hb8 == io_inputs_1 ? 7'h64 : _GEN_2487; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2489 = 10'hb9 == io_inputs_1 ? 7'h64 : _GEN_2488; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2490 = 10'hba == io_inputs_1 ? 7'h64 : _GEN_2489; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2491 = 10'hbb == io_inputs_1 ? 7'h64 : _GEN_2490; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2492 = 10'hbc == io_inputs_1 ? 7'h64 : _GEN_2491; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2493 = 10'hbd == io_inputs_1 ? 7'h64 : _GEN_2492; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2494 = 10'hbe == io_inputs_1 ? 7'h64 : _GEN_2493; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2495 = 10'hbf == io_inputs_1 ? 7'h64 : _GEN_2494; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2496 = 10'hc0 == io_inputs_1 ? 7'h64 : _GEN_2495; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2497 = 10'hc1 == io_inputs_1 ? 7'h64 : _GEN_2496; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2498 = 10'hc2 == io_inputs_1 ? 7'h64 : _GEN_2497; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2499 = 10'hc3 == io_inputs_1 ? 7'h64 : _GEN_2498; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2500 = 10'hc4 == io_inputs_1 ? 7'h64 : _GEN_2499; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2501 = 10'hc5 == io_inputs_1 ? 7'h64 : _GEN_2500; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2502 = 10'hc6 == io_inputs_1 ? 7'h64 : _GEN_2501; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2503 = 10'hc7 == io_inputs_1 ? 7'h64 : _GEN_2502; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2504 = 10'hc8 == io_inputs_1 ? 7'h64 : _GEN_2503; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2505 = 10'hc9 == io_inputs_1 ? 7'h63 : _GEN_2504; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2506 = 10'hca == io_inputs_1 ? 7'h62 : _GEN_2505; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2507 = 10'hcb == io_inputs_1 ? 7'h61 : _GEN_2506; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2508 = 10'hcc == io_inputs_1 ? 7'h60 : _GEN_2507; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2509 = 10'hcd == io_inputs_1 ? 7'h5f : _GEN_2508; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2510 = 10'hce == io_inputs_1 ? 7'h5e : _GEN_2509; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2511 = 10'hcf == io_inputs_1 ? 7'h5d : _GEN_2510; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2512 = 10'hd0 == io_inputs_1 ? 7'h5c : _GEN_2511; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2513 = 10'hd1 == io_inputs_1 ? 7'h5b : _GEN_2512; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2514 = 10'hd2 == io_inputs_1 ? 7'h5a : _GEN_2513; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2515 = 10'hd3 == io_inputs_1 ? 7'h59 : _GEN_2514; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2516 = 10'hd4 == io_inputs_1 ? 7'h58 : _GEN_2515; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2517 = 10'hd5 == io_inputs_1 ? 7'h57 : _GEN_2516; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2518 = 10'hd6 == io_inputs_1 ? 7'h56 : _GEN_2517; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2519 = 10'hd7 == io_inputs_1 ? 7'h55 : _GEN_2518; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2520 = 10'hd8 == io_inputs_1 ? 7'h54 : _GEN_2519; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2521 = 10'hd9 == io_inputs_1 ? 7'h53 : _GEN_2520; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2522 = 10'hda == io_inputs_1 ? 7'h52 : _GEN_2521; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2523 = 10'hdb == io_inputs_1 ? 7'h51 : _GEN_2522; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2524 = 10'hdc == io_inputs_1 ? 7'h50 : _GEN_2523; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2525 = 10'hdd == io_inputs_1 ? 7'h4f : _GEN_2524; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2526 = 10'hde == io_inputs_1 ? 7'h4e : _GEN_2525; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2527 = 10'hdf == io_inputs_1 ? 7'h4d : _GEN_2526; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2528 = 10'he0 == io_inputs_1 ? 7'h4c : _GEN_2527; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2529 = 10'he1 == io_inputs_1 ? 7'h4b : _GEN_2528; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2530 = 10'he2 == io_inputs_1 ? 7'h4a : _GEN_2529; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2531 = 10'he3 == io_inputs_1 ? 7'h49 : _GEN_2530; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2532 = 10'he4 == io_inputs_1 ? 7'h48 : _GEN_2531; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2533 = 10'he5 == io_inputs_1 ? 7'h47 : _GEN_2532; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2534 = 10'he6 == io_inputs_1 ? 7'h46 : _GEN_2533; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2535 = 10'he7 == io_inputs_1 ? 7'h45 : _GEN_2534; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2536 = 10'he8 == io_inputs_1 ? 7'h44 : _GEN_2535; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2537 = 10'he9 == io_inputs_1 ? 7'h43 : _GEN_2536; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2538 = 10'hea == io_inputs_1 ? 7'h42 : _GEN_2537; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2539 = 10'heb == io_inputs_1 ? 7'h41 : _GEN_2538; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2540 = 10'hec == io_inputs_1 ? 7'h40 : _GEN_2539; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2541 = 10'hed == io_inputs_1 ? 7'h3f : _GEN_2540; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2542 = 10'hee == io_inputs_1 ? 7'h3e : _GEN_2541; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2543 = 10'hef == io_inputs_1 ? 7'h3d : _GEN_2542; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2544 = 10'hf0 == io_inputs_1 ? 7'h3c : _GEN_2543; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2545 = 10'hf1 == io_inputs_1 ? 7'h3b : _GEN_2544; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2546 = 10'hf2 == io_inputs_1 ? 7'h3a : _GEN_2545; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2547 = 10'hf3 == io_inputs_1 ? 7'h39 : _GEN_2546; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2548 = 10'hf4 == io_inputs_1 ? 7'h38 : _GEN_2547; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2549 = 10'hf5 == io_inputs_1 ? 7'h37 : _GEN_2548; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2550 = 10'hf6 == io_inputs_1 ? 7'h36 : _GEN_2549; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2551 = 10'hf7 == io_inputs_1 ? 7'h35 : _GEN_2550; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2552 = 10'hf8 == io_inputs_1 ? 7'h34 : _GEN_2551; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2553 = 10'hf9 == io_inputs_1 ? 7'h33 : _GEN_2552; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2554 = 10'hfa == io_inputs_1 ? 7'h32 : _GEN_2553; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2555 = 10'hfb == io_inputs_1 ? 7'h31 : _GEN_2554; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2556 = 10'hfc == io_inputs_1 ? 7'h30 : _GEN_2555; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2557 = 10'hfd == io_inputs_1 ? 7'h2f : _GEN_2556; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2558 = 10'hfe == io_inputs_1 ? 7'h2e : _GEN_2557; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2559 = 10'hff == io_inputs_1 ? 7'h2d : _GEN_2558; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2560 = 10'h100 == io_inputs_1 ? 7'h2c : _GEN_2559; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2561 = 10'h101 == io_inputs_1 ? 7'h2b : _GEN_2560; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2562 = 10'h102 == io_inputs_1 ? 7'h2a : _GEN_2561; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2563 = 10'h103 == io_inputs_1 ? 7'h29 : _GEN_2562; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2564 = 10'h104 == io_inputs_1 ? 7'h28 : _GEN_2563; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2565 = 10'h105 == io_inputs_1 ? 7'h27 : _GEN_2564; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2566 = 10'h106 == io_inputs_1 ? 7'h26 : _GEN_2565; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2567 = 10'h107 == io_inputs_1 ? 7'h25 : _GEN_2566; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2568 = 10'h108 == io_inputs_1 ? 7'h24 : _GEN_2567; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2569 = 10'h109 == io_inputs_1 ? 7'h23 : _GEN_2568; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2570 = 10'h10a == io_inputs_1 ? 7'h22 : _GEN_2569; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2571 = 10'h10b == io_inputs_1 ? 7'h21 : _GEN_2570; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2572 = 10'h10c == io_inputs_1 ? 7'h20 : _GEN_2571; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2573 = 10'h10d == io_inputs_1 ? 7'h1f : _GEN_2572; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2574 = 10'h10e == io_inputs_1 ? 7'h1e : _GEN_2573; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2575 = 10'h10f == io_inputs_1 ? 7'h1d : _GEN_2574; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2576 = 10'h110 == io_inputs_1 ? 7'h1c : _GEN_2575; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2577 = 10'h111 == io_inputs_1 ? 7'h1b : _GEN_2576; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2578 = 10'h112 == io_inputs_1 ? 7'h1a : _GEN_2577; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2579 = 10'h113 == io_inputs_1 ? 7'h19 : _GEN_2578; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2580 = 10'h114 == io_inputs_1 ? 7'h18 : _GEN_2579; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2581 = 10'h115 == io_inputs_1 ? 7'h17 : _GEN_2580; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2582 = 10'h116 == io_inputs_1 ? 7'h16 : _GEN_2581; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2583 = 10'h117 == io_inputs_1 ? 7'h15 : _GEN_2582; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2584 = 10'h118 == io_inputs_1 ? 7'h14 : _GEN_2583; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2585 = 10'h119 == io_inputs_1 ? 7'h13 : _GEN_2584; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2586 = 10'h11a == io_inputs_1 ? 7'h12 : _GEN_2585; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2587 = 10'h11b == io_inputs_1 ? 7'h11 : _GEN_2586; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2588 = 10'h11c == io_inputs_1 ? 7'h10 : _GEN_2587; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2589 = 10'h11d == io_inputs_1 ? 7'hf : _GEN_2588; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2590 = 10'h11e == io_inputs_1 ? 7'he : _GEN_2589; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2591 = 10'h11f == io_inputs_1 ? 7'hd : _GEN_2590; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2592 = 10'h120 == io_inputs_1 ? 7'hc : _GEN_2591; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2593 = 10'h121 == io_inputs_1 ? 7'hb : _GEN_2592; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2594 = 10'h122 == io_inputs_1 ? 7'ha : _GEN_2593; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2595 = 10'h123 == io_inputs_1 ? 7'h9 : _GEN_2594; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2596 = 10'h124 == io_inputs_1 ? 7'h8 : _GEN_2595; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2597 = 10'h125 == io_inputs_1 ? 7'h7 : _GEN_2596; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2598 = 10'h126 == io_inputs_1 ? 7'h6 : _GEN_2597; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2599 = 10'h127 == io_inputs_1 ? 7'h5 : _GEN_2598; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2600 = 10'h128 == io_inputs_1 ? 7'h4 : _GEN_2599; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2601 = 10'h129 == io_inputs_1 ? 7'h3 : _GEN_2600; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2602 = 10'h12a == io_inputs_1 ? 7'h2 : _GEN_2601; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2603 = 10'h12b == io_inputs_1 ? 7'h1 : _GEN_2602; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2604 = 10'h12c == io_inputs_1 ? 7'h0 : _GEN_2603; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2605 = 10'h12d == io_inputs_1 ? 7'h0 : _GEN_2604; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2606 = 10'h12e == io_inputs_1 ? 7'h0 : _GEN_2605; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2607 = 10'h12f == io_inputs_1 ? 7'h0 : _GEN_2606; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2608 = 10'h130 == io_inputs_1 ? 7'h0 : _GEN_2607; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2609 = 10'h131 == io_inputs_1 ? 7'h0 : _GEN_2608; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2610 = 10'h132 == io_inputs_1 ? 7'h0 : _GEN_2609; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2611 = 10'h133 == io_inputs_1 ? 7'h0 : _GEN_2610; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2612 = 10'h134 == io_inputs_1 ? 7'h0 : _GEN_2611; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2613 = 10'h135 == io_inputs_1 ? 7'h0 : _GEN_2612; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2614 = 10'h136 == io_inputs_1 ? 7'h0 : _GEN_2613; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2615 = 10'h137 == io_inputs_1 ? 7'h0 : _GEN_2614; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2616 = 10'h138 == io_inputs_1 ? 7'h0 : _GEN_2615; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2617 = 10'h139 == io_inputs_1 ? 7'h0 : _GEN_2616; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2618 = 10'h13a == io_inputs_1 ? 7'h0 : _GEN_2617; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2619 = 10'h13b == io_inputs_1 ? 7'h0 : _GEN_2618; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2620 = 10'h13c == io_inputs_1 ? 7'h0 : _GEN_2619; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2621 = 10'h13d == io_inputs_1 ? 7'h0 : _GEN_2620; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2622 = 10'h13e == io_inputs_1 ? 7'h0 : _GEN_2621; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2623 = 10'h13f == io_inputs_1 ? 7'h0 : _GEN_2622; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2624 = 10'h140 == io_inputs_1 ? 7'h0 : _GEN_2623; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2625 = 10'h141 == io_inputs_1 ? 7'h0 : _GEN_2624; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2626 = 10'h142 == io_inputs_1 ? 7'h0 : _GEN_2625; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2627 = 10'h143 == io_inputs_1 ? 7'h0 : _GEN_2626; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2628 = 10'h144 == io_inputs_1 ? 7'h0 : _GEN_2627; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2629 = 10'h145 == io_inputs_1 ? 7'h0 : _GEN_2628; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2630 = 10'h146 == io_inputs_1 ? 7'h0 : _GEN_2629; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2631 = 10'h147 == io_inputs_1 ? 7'h0 : _GEN_2630; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2632 = 10'h148 == io_inputs_1 ? 7'h0 : _GEN_2631; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2633 = 10'h149 == io_inputs_1 ? 7'h0 : _GEN_2632; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2634 = 10'h14a == io_inputs_1 ? 7'h0 : _GEN_2633; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2635 = 10'h14b == io_inputs_1 ? 7'h0 : _GEN_2634; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2636 = 10'h14c == io_inputs_1 ? 7'h0 : _GEN_2635; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2637 = 10'h14d == io_inputs_1 ? 7'h0 : _GEN_2636; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2638 = 10'h14e == io_inputs_1 ? 7'h0 : _GEN_2637; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2639 = 10'h14f == io_inputs_1 ? 7'h0 : _GEN_2638; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2640 = 10'h150 == io_inputs_1 ? 7'h0 : _GEN_2639; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2641 = 10'h151 == io_inputs_1 ? 7'h0 : _GEN_2640; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2642 = 10'h152 == io_inputs_1 ? 7'h0 : _GEN_2641; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2643 = 10'h153 == io_inputs_1 ? 7'h0 : _GEN_2642; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2644 = 10'h154 == io_inputs_1 ? 7'h0 : _GEN_2643; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2645 = 10'h155 == io_inputs_1 ? 7'h0 : _GEN_2644; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2646 = 10'h156 == io_inputs_1 ? 7'h0 : _GEN_2645; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2647 = 10'h157 == io_inputs_1 ? 7'h0 : _GEN_2646; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2648 = 10'h158 == io_inputs_1 ? 7'h0 : _GEN_2647; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2649 = 10'h159 == io_inputs_1 ? 7'h0 : _GEN_2648; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2650 = 10'h15a == io_inputs_1 ? 7'h0 : _GEN_2649; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2651 = 10'h15b == io_inputs_1 ? 7'h0 : _GEN_2650; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2652 = 10'h15c == io_inputs_1 ? 7'h0 : _GEN_2651; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2653 = 10'h15d == io_inputs_1 ? 7'h0 : _GEN_2652; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2654 = 10'h15e == io_inputs_1 ? 7'h0 : _GEN_2653; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2655 = 10'h15f == io_inputs_1 ? 7'h0 : _GEN_2654; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2656 = 10'h160 == io_inputs_1 ? 7'h0 : _GEN_2655; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2657 = 10'h161 == io_inputs_1 ? 7'h0 : _GEN_2656; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2658 = 10'h162 == io_inputs_1 ? 7'h0 : _GEN_2657; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2659 = 10'h163 == io_inputs_1 ? 7'h0 : _GEN_2658; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2660 = 10'h164 == io_inputs_1 ? 7'h0 : _GEN_2659; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2661 = 10'h165 == io_inputs_1 ? 7'h0 : _GEN_2660; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2662 = 10'h166 == io_inputs_1 ? 7'h0 : _GEN_2661; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2663 = 10'h167 == io_inputs_1 ? 7'h0 : _GEN_2662; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2664 = 10'h168 == io_inputs_1 ? 7'h0 : _GEN_2663; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2665 = 10'h169 == io_inputs_1 ? 7'h0 : _GEN_2664; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2666 = 10'h16a == io_inputs_1 ? 7'h0 : _GEN_2665; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2667 = 10'h16b == io_inputs_1 ? 7'h0 : _GEN_2666; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2668 = 10'h16c == io_inputs_1 ? 7'h0 : _GEN_2667; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2669 = 10'h16d == io_inputs_1 ? 7'h0 : _GEN_2668; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2670 = 10'h16e == io_inputs_1 ? 7'h0 : _GEN_2669; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2671 = 10'h16f == io_inputs_1 ? 7'h0 : _GEN_2670; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2672 = 10'h170 == io_inputs_1 ? 7'h0 : _GEN_2671; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2673 = 10'h171 == io_inputs_1 ? 7'h0 : _GEN_2672; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2674 = 10'h172 == io_inputs_1 ? 7'h0 : _GEN_2673; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2675 = 10'h173 == io_inputs_1 ? 7'h0 : _GEN_2674; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2676 = 10'h174 == io_inputs_1 ? 7'h0 : _GEN_2675; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2677 = 10'h175 == io_inputs_1 ? 7'h0 : _GEN_2676; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2678 = 10'h176 == io_inputs_1 ? 7'h0 : _GEN_2677; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2679 = 10'h177 == io_inputs_1 ? 7'h0 : _GEN_2678; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2680 = 10'h178 == io_inputs_1 ? 7'h0 : _GEN_2679; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2681 = 10'h179 == io_inputs_1 ? 7'h0 : _GEN_2680; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2682 = 10'h17a == io_inputs_1 ? 7'h0 : _GEN_2681; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2683 = 10'h17b == io_inputs_1 ? 7'h0 : _GEN_2682; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2684 = 10'h17c == io_inputs_1 ? 7'h0 : _GEN_2683; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2685 = 10'h17d == io_inputs_1 ? 7'h0 : _GEN_2684; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2686 = 10'h17e == io_inputs_1 ? 7'h0 : _GEN_2685; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2687 = 10'h17f == io_inputs_1 ? 7'h0 : _GEN_2686; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2688 = 10'h180 == io_inputs_1 ? 7'h0 : _GEN_2687; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2689 = 10'h181 == io_inputs_1 ? 7'h0 : _GEN_2688; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2690 = 10'h182 == io_inputs_1 ? 7'h0 : _GEN_2689; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2691 = 10'h183 == io_inputs_1 ? 7'h0 : _GEN_2690; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2692 = 10'h184 == io_inputs_1 ? 7'h0 : _GEN_2691; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2693 = 10'h185 == io_inputs_1 ? 7'h0 : _GEN_2692; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2694 = 10'h186 == io_inputs_1 ? 7'h0 : _GEN_2693; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2695 = 10'h187 == io_inputs_1 ? 7'h0 : _GEN_2694; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2696 = 10'h188 == io_inputs_1 ? 7'h0 : _GEN_2695; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2697 = 10'h189 == io_inputs_1 ? 7'h0 : _GEN_2696; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2698 = 10'h18a == io_inputs_1 ? 7'h0 : _GEN_2697; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2699 = 10'h18b == io_inputs_1 ? 7'h0 : _GEN_2698; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2700 = 10'h18c == io_inputs_1 ? 7'h0 : _GEN_2699; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2701 = 10'h18d == io_inputs_1 ? 7'h0 : _GEN_2700; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2702 = 10'h18e == io_inputs_1 ? 7'h0 : _GEN_2701; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2703 = 10'h18f == io_inputs_1 ? 7'h0 : _GEN_2702; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2704 = 10'h190 == io_inputs_1 ? 7'h0 : _GEN_2703; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2705 = 10'h191 == io_inputs_1 ? 7'h0 : _GEN_2704; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2706 = 10'h192 == io_inputs_1 ? 7'h0 : _GEN_2705; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2707 = 10'h193 == io_inputs_1 ? 7'h0 : _GEN_2706; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2708 = 10'h194 == io_inputs_1 ? 7'h0 : _GEN_2707; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2709 = 10'h195 == io_inputs_1 ? 7'h0 : _GEN_2708; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2710 = 10'h196 == io_inputs_1 ? 7'h0 : _GEN_2709; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2711 = 10'h197 == io_inputs_1 ? 7'h0 : _GEN_2710; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2712 = 10'h198 == io_inputs_1 ? 7'h0 : _GEN_2711; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2713 = 10'h199 == io_inputs_1 ? 7'h0 : _GEN_2712; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2714 = 10'h19a == io_inputs_1 ? 7'h0 : _GEN_2713; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2715 = 10'h19b == io_inputs_1 ? 7'h0 : _GEN_2714; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2716 = 10'h19c == io_inputs_1 ? 7'h0 : _GEN_2715; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2717 = 10'h19d == io_inputs_1 ? 7'h0 : _GEN_2716; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2718 = 10'h19e == io_inputs_1 ? 7'h0 : _GEN_2717; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2719 = 10'h19f == io_inputs_1 ? 7'h0 : _GEN_2718; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2720 = 10'h1a0 == io_inputs_1 ? 7'h0 : _GEN_2719; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2721 = 10'h1a1 == io_inputs_1 ? 7'h0 : _GEN_2720; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2722 = 10'h1a2 == io_inputs_1 ? 7'h0 : _GEN_2721; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2723 = 10'h1a3 == io_inputs_1 ? 7'h0 : _GEN_2722; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2724 = 10'h1a4 == io_inputs_1 ? 7'h0 : _GEN_2723; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2725 = 10'h1a5 == io_inputs_1 ? 7'h0 : _GEN_2724; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2726 = 10'h1a6 == io_inputs_1 ? 7'h0 : _GEN_2725; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2727 = 10'h1a7 == io_inputs_1 ? 7'h0 : _GEN_2726; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2728 = 10'h1a8 == io_inputs_1 ? 7'h0 : _GEN_2727; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2729 = 10'h1a9 == io_inputs_1 ? 7'h0 : _GEN_2728; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2730 = 10'h1aa == io_inputs_1 ? 7'h0 : _GEN_2729; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2731 = 10'h1ab == io_inputs_1 ? 7'h0 : _GEN_2730; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2732 = 10'h1ac == io_inputs_1 ? 7'h0 : _GEN_2731; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2733 = 10'h1ad == io_inputs_1 ? 7'h0 : _GEN_2732; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2734 = 10'h1ae == io_inputs_1 ? 7'h0 : _GEN_2733; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2735 = 10'h1af == io_inputs_1 ? 7'h0 : _GEN_2734; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2736 = 10'h1b0 == io_inputs_1 ? 7'h0 : _GEN_2735; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2737 = 10'h1b1 == io_inputs_1 ? 7'h0 : _GEN_2736; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2738 = 10'h1b2 == io_inputs_1 ? 7'h0 : _GEN_2737; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2739 = 10'h1b3 == io_inputs_1 ? 7'h0 : _GEN_2738; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2740 = 10'h1b4 == io_inputs_1 ? 7'h0 : _GEN_2739; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2741 = 10'h1b5 == io_inputs_1 ? 7'h0 : _GEN_2740; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2742 = 10'h1b6 == io_inputs_1 ? 7'h0 : _GEN_2741; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2743 = 10'h1b7 == io_inputs_1 ? 7'h0 : _GEN_2742; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2744 = 10'h1b8 == io_inputs_1 ? 7'h0 : _GEN_2743; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2745 = 10'h1b9 == io_inputs_1 ? 7'h0 : _GEN_2744; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2746 = 10'h1ba == io_inputs_1 ? 7'h0 : _GEN_2745; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2747 = 10'h1bb == io_inputs_1 ? 7'h0 : _GEN_2746; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2748 = 10'h1bc == io_inputs_1 ? 7'h0 : _GEN_2747; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2749 = 10'h1bd == io_inputs_1 ? 7'h0 : _GEN_2748; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2750 = 10'h1be == io_inputs_1 ? 7'h0 : _GEN_2749; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2751 = 10'h1bf == io_inputs_1 ? 7'h0 : _GEN_2750; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2752 = 10'h1c0 == io_inputs_1 ? 7'h0 : _GEN_2751; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2753 = 10'h1c1 == io_inputs_1 ? 7'h0 : _GEN_2752; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2754 = 10'h1c2 == io_inputs_1 ? 7'h0 : _GEN_2753; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2755 = 10'h1c3 == io_inputs_1 ? 7'h0 : _GEN_2754; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2756 = 10'h1c4 == io_inputs_1 ? 7'h0 : _GEN_2755; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2757 = 10'h1c5 == io_inputs_1 ? 7'h0 : _GEN_2756; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2758 = 10'h1c6 == io_inputs_1 ? 7'h0 : _GEN_2757; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2759 = 10'h1c7 == io_inputs_1 ? 7'h0 : _GEN_2758; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2760 = 10'h1c8 == io_inputs_1 ? 7'h0 : _GEN_2759; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2761 = 10'h1c9 == io_inputs_1 ? 7'h0 : _GEN_2760; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2762 = 10'h1ca == io_inputs_1 ? 7'h0 : _GEN_2761; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2763 = 10'h1cb == io_inputs_1 ? 7'h0 : _GEN_2762; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2764 = 10'h1cc == io_inputs_1 ? 7'h0 : _GEN_2763; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2765 = 10'h1cd == io_inputs_1 ? 7'h0 : _GEN_2764; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2766 = 10'h1ce == io_inputs_1 ? 7'h0 : _GEN_2765; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2767 = 10'h1cf == io_inputs_1 ? 7'h0 : _GEN_2766; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2768 = 10'h1d0 == io_inputs_1 ? 7'h0 : _GEN_2767; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2769 = 10'h1d1 == io_inputs_1 ? 7'h0 : _GEN_2768; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2770 = 10'h1d2 == io_inputs_1 ? 7'h0 : _GEN_2769; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2771 = 10'h1d3 == io_inputs_1 ? 7'h0 : _GEN_2770; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2772 = 10'h1d4 == io_inputs_1 ? 7'h0 : _GEN_2771; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2773 = 10'h1d5 == io_inputs_1 ? 7'h0 : _GEN_2772; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2774 = 10'h1d6 == io_inputs_1 ? 7'h0 : _GEN_2773; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2775 = 10'h1d7 == io_inputs_1 ? 7'h0 : _GEN_2774; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2776 = 10'h1d8 == io_inputs_1 ? 7'h0 : _GEN_2775; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2777 = 10'h1d9 == io_inputs_1 ? 7'h0 : _GEN_2776; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2778 = 10'h1da == io_inputs_1 ? 7'h0 : _GEN_2777; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2779 = 10'h1db == io_inputs_1 ? 7'h0 : _GEN_2778; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2780 = 10'h1dc == io_inputs_1 ? 7'h0 : _GEN_2779; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2781 = 10'h1dd == io_inputs_1 ? 7'h0 : _GEN_2780; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2782 = 10'h1de == io_inputs_1 ? 7'h0 : _GEN_2781; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2783 = 10'h1df == io_inputs_1 ? 7'h0 : _GEN_2782; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2784 = 10'h1e0 == io_inputs_1 ? 7'h0 : _GEN_2783; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2785 = 10'h1e1 == io_inputs_1 ? 7'h0 : _GEN_2784; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2786 = 10'h1e2 == io_inputs_1 ? 7'h0 : _GEN_2785; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2787 = 10'h1e3 == io_inputs_1 ? 7'h0 : _GEN_2786; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2788 = 10'h1e4 == io_inputs_1 ? 7'h0 : _GEN_2787; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2789 = 10'h1e5 == io_inputs_1 ? 7'h0 : _GEN_2788; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2790 = 10'h1e6 == io_inputs_1 ? 7'h0 : _GEN_2789; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2791 = 10'h1e7 == io_inputs_1 ? 7'h0 : _GEN_2790; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2792 = 10'h1e8 == io_inputs_1 ? 7'h0 : _GEN_2791; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2793 = 10'h1e9 == io_inputs_1 ? 7'h0 : _GEN_2792; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2794 = 10'h1ea == io_inputs_1 ? 7'h0 : _GEN_2793; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2795 = 10'h1eb == io_inputs_1 ? 7'h0 : _GEN_2794; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2796 = 10'h1ec == io_inputs_1 ? 7'h0 : _GEN_2795; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2797 = 10'h1ed == io_inputs_1 ? 7'h0 : _GEN_2796; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2798 = 10'h1ee == io_inputs_1 ? 7'h0 : _GEN_2797; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2799 = 10'h1ef == io_inputs_1 ? 7'h0 : _GEN_2798; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2800 = 10'h1f0 == io_inputs_1 ? 7'h0 : _GEN_2799; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2801 = 10'h1f1 == io_inputs_1 ? 7'h0 : _GEN_2800; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2802 = 10'h1f2 == io_inputs_1 ? 7'h0 : _GEN_2801; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2803 = 10'h1f3 == io_inputs_1 ? 7'h0 : _GEN_2802; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2804 = 10'h1f4 == io_inputs_1 ? 7'h0 : _GEN_2803; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2805 = 10'h1f5 == io_inputs_1 ? 7'h0 : _GEN_2804; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2806 = 10'h1f6 == io_inputs_1 ? 7'h0 : _GEN_2805; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2807 = 10'h1f7 == io_inputs_1 ? 7'h0 : _GEN_2806; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2808 = 10'h1f8 == io_inputs_1 ? 7'h0 : _GEN_2807; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2809 = 10'h1f9 == io_inputs_1 ? 7'h0 : _GEN_2808; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2810 = 10'h1fa == io_inputs_1 ? 7'h0 : _GEN_2809; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2811 = 10'h1fb == io_inputs_1 ? 7'h0 : _GEN_2810; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2812 = 10'h1fc == io_inputs_1 ? 7'h0 : _GEN_2811; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2813 = 10'h1fd == io_inputs_1 ? 7'h0 : _GEN_2812; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2814 = 10'h1fe == io_inputs_1 ? 7'h0 : _GEN_2813; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2815 = 10'h1ff == io_inputs_1 ? 7'h0 : _GEN_2814; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2816 = 10'h200 == io_inputs_1 ? 7'h0 : _GEN_2815; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2817 = 10'h201 == io_inputs_1 ? 7'h0 : _GEN_2816; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2818 = 10'h202 == io_inputs_1 ? 7'h0 : _GEN_2817; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2819 = 10'h203 == io_inputs_1 ? 7'h0 : _GEN_2818; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2820 = 10'h204 == io_inputs_1 ? 7'h0 : _GEN_2819; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2821 = 10'h205 == io_inputs_1 ? 7'h0 : _GEN_2820; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2822 = 10'h206 == io_inputs_1 ? 7'h0 : _GEN_2821; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2823 = 10'h207 == io_inputs_1 ? 7'h0 : _GEN_2822; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2824 = 10'h208 == io_inputs_1 ? 7'h0 : _GEN_2823; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2825 = 10'h209 == io_inputs_1 ? 7'h0 : _GEN_2824; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2826 = 10'h20a == io_inputs_1 ? 7'h0 : _GEN_2825; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2827 = 10'h20b == io_inputs_1 ? 7'h0 : _GEN_2826; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2828 = 10'h20c == io_inputs_1 ? 7'h0 : _GEN_2827; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2829 = 10'h20d == io_inputs_1 ? 7'h0 : _GEN_2828; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2830 = 10'h20e == io_inputs_1 ? 7'h0 : _GEN_2829; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2831 = 10'h20f == io_inputs_1 ? 7'h0 : _GEN_2830; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2832 = 10'h210 == io_inputs_1 ? 7'h0 : _GEN_2831; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2833 = 10'h211 == io_inputs_1 ? 7'h0 : _GEN_2832; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2834 = 10'h212 == io_inputs_1 ? 7'h0 : _GEN_2833; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2835 = 10'h213 == io_inputs_1 ? 7'h0 : _GEN_2834; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2836 = 10'h214 == io_inputs_1 ? 7'h0 : _GEN_2835; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2837 = 10'h215 == io_inputs_1 ? 7'h0 : _GEN_2836; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2838 = 10'h216 == io_inputs_1 ? 7'h0 : _GEN_2837; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2839 = 10'h217 == io_inputs_1 ? 7'h0 : _GEN_2838; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2840 = 10'h218 == io_inputs_1 ? 7'h0 : _GEN_2839; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2841 = 10'h219 == io_inputs_1 ? 7'h0 : _GEN_2840; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2842 = 10'h21a == io_inputs_1 ? 7'h0 : _GEN_2841; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2843 = 10'h21b == io_inputs_1 ? 7'h0 : _GEN_2842; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2844 = 10'h21c == io_inputs_1 ? 7'h0 : _GEN_2843; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2845 = 10'h21d == io_inputs_1 ? 7'h0 : _GEN_2844; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2846 = 10'h21e == io_inputs_1 ? 7'h0 : _GEN_2845; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2847 = 10'h21f == io_inputs_1 ? 7'h0 : _GEN_2846; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2848 = 10'h220 == io_inputs_1 ? 7'h0 : _GEN_2847; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2849 = 10'h221 == io_inputs_1 ? 7'h0 : _GEN_2848; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2850 = 10'h222 == io_inputs_1 ? 7'h0 : _GEN_2849; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2851 = 10'h223 == io_inputs_1 ? 7'h0 : _GEN_2850; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2852 = 10'h224 == io_inputs_1 ? 7'h0 : _GEN_2851; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2853 = 10'h225 == io_inputs_1 ? 7'h0 : _GEN_2852; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2854 = 10'h226 == io_inputs_1 ? 7'h0 : _GEN_2853; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2855 = 10'h227 == io_inputs_1 ? 7'h0 : _GEN_2854; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2856 = 10'h228 == io_inputs_1 ? 7'h0 : _GEN_2855; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2857 = 10'h229 == io_inputs_1 ? 7'h0 : _GEN_2856; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2858 = 10'h22a == io_inputs_1 ? 7'h0 : _GEN_2857; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2859 = 10'h22b == io_inputs_1 ? 7'h0 : _GEN_2858; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2860 = 10'h22c == io_inputs_1 ? 7'h0 : _GEN_2859; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2861 = 10'h22d == io_inputs_1 ? 7'h0 : _GEN_2860; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2862 = 10'h22e == io_inputs_1 ? 7'h0 : _GEN_2861; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2863 = 10'h22f == io_inputs_1 ? 7'h0 : _GEN_2862; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2864 = 10'h230 == io_inputs_1 ? 7'h0 : _GEN_2863; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2865 = 10'h231 == io_inputs_1 ? 7'h0 : _GEN_2864; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2866 = 10'h232 == io_inputs_1 ? 7'h0 : _GEN_2865; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2867 = 10'h233 == io_inputs_1 ? 7'h0 : _GEN_2866; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2868 = 10'h234 == io_inputs_1 ? 7'h0 : _GEN_2867; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2869 = 10'h235 == io_inputs_1 ? 7'h0 : _GEN_2868; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2870 = 10'h236 == io_inputs_1 ? 7'h0 : _GEN_2869; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2871 = 10'h237 == io_inputs_1 ? 7'h0 : _GEN_2870; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2872 = 10'h238 == io_inputs_1 ? 7'h0 : _GEN_2871; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2873 = 10'h239 == io_inputs_1 ? 7'h0 : _GEN_2872; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2874 = 10'h23a == io_inputs_1 ? 7'h0 : _GEN_2873; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2875 = 10'h23b == io_inputs_1 ? 7'h0 : _GEN_2874; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2876 = 10'h23c == io_inputs_1 ? 7'h0 : _GEN_2875; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2877 = 10'h23d == io_inputs_1 ? 7'h0 : _GEN_2876; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2878 = 10'h23e == io_inputs_1 ? 7'h0 : _GEN_2877; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2879 = 10'h23f == io_inputs_1 ? 7'h0 : _GEN_2878; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2880 = 10'h240 == io_inputs_1 ? 7'h0 : _GEN_2879; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2881 = 10'h241 == io_inputs_1 ? 7'h0 : _GEN_2880; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2882 = 10'h242 == io_inputs_1 ? 7'h0 : _GEN_2881; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2883 = 10'h243 == io_inputs_1 ? 7'h0 : _GEN_2882; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2884 = 10'h244 == io_inputs_1 ? 7'h0 : _GEN_2883; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2885 = 10'h245 == io_inputs_1 ? 7'h0 : _GEN_2884; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2886 = 10'h246 == io_inputs_1 ? 7'h0 : _GEN_2885; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2887 = 10'h247 == io_inputs_1 ? 7'h0 : _GEN_2886; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2888 = 10'h248 == io_inputs_1 ? 7'h0 : _GEN_2887; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2889 = 10'h249 == io_inputs_1 ? 7'h0 : _GEN_2888; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2890 = 10'h24a == io_inputs_1 ? 7'h0 : _GEN_2889; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2891 = 10'h24b == io_inputs_1 ? 7'h0 : _GEN_2890; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2892 = 10'h24c == io_inputs_1 ? 7'h0 : _GEN_2891; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2893 = 10'h24d == io_inputs_1 ? 7'h0 : _GEN_2892; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2894 = 10'h24e == io_inputs_1 ? 7'h0 : _GEN_2893; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2895 = 10'h24f == io_inputs_1 ? 7'h0 : _GEN_2894; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2896 = 10'h250 == io_inputs_1 ? 7'h0 : _GEN_2895; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2897 = 10'h251 == io_inputs_1 ? 7'h0 : _GEN_2896; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2898 = 10'h252 == io_inputs_1 ? 7'h0 : _GEN_2897; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2899 = 10'h253 == io_inputs_1 ? 7'h0 : _GEN_2898; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2900 = 10'h254 == io_inputs_1 ? 7'h0 : _GEN_2899; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2901 = 10'h255 == io_inputs_1 ? 7'h0 : _GEN_2900; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2902 = 10'h256 == io_inputs_1 ? 7'h0 : _GEN_2901; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2903 = 10'h257 == io_inputs_1 ? 7'h0 : _GEN_2902; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2904 = 10'h258 == io_inputs_1 ? 7'h0 : _GEN_2903; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2905 = 10'h259 == io_inputs_1 ? 7'h0 : _GEN_2904; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2906 = 10'h25a == io_inputs_1 ? 7'h0 : _GEN_2905; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2907 = 10'h25b == io_inputs_1 ? 7'h0 : _GEN_2906; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2908 = 10'h25c == io_inputs_1 ? 7'h0 : _GEN_2907; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2909 = 10'h25d == io_inputs_1 ? 7'h0 : _GEN_2908; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2910 = 10'h25e == io_inputs_1 ? 7'h0 : _GEN_2909; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2911 = 10'h25f == io_inputs_1 ? 7'h0 : _GEN_2910; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2912 = 10'h260 == io_inputs_1 ? 7'h0 : _GEN_2911; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2913 = 10'h261 == io_inputs_1 ? 7'h0 : _GEN_2912; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2914 = 10'h262 == io_inputs_1 ? 7'h0 : _GEN_2913; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2915 = 10'h263 == io_inputs_1 ? 7'h0 : _GEN_2914; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2916 = 10'h264 == io_inputs_1 ? 7'h0 : _GEN_2915; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2917 = 10'h265 == io_inputs_1 ? 7'h0 : _GEN_2916; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2918 = 10'h266 == io_inputs_1 ? 7'h0 : _GEN_2917; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2919 = 10'h267 == io_inputs_1 ? 7'h0 : _GEN_2918; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2920 = 10'h268 == io_inputs_1 ? 7'h0 : _GEN_2919; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2921 = 10'h269 == io_inputs_1 ? 7'h0 : _GEN_2920; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2922 = 10'h26a == io_inputs_1 ? 7'h0 : _GEN_2921; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2923 = 10'h26b == io_inputs_1 ? 7'h0 : _GEN_2922; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2924 = 10'h26c == io_inputs_1 ? 7'h0 : _GEN_2923; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2925 = 10'h26d == io_inputs_1 ? 7'h0 : _GEN_2924; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2926 = 10'h26e == io_inputs_1 ? 7'h0 : _GEN_2925; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2927 = 10'h26f == io_inputs_1 ? 7'h0 : _GEN_2926; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2928 = 10'h270 == io_inputs_1 ? 7'h0 : _GEN_2927; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2929 = 10'h271 == io_inputs_1 ? 7'h0 : _GEN_2928; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2930 = 10'h272 == io_inputs_1 ? 7'h0 : _GEN_2929; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2931 = 10'h273 == io_inputs_1 ? 7'h0 : _GEN_2930; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2932 = 10'h274 == io_inputs_1 ? 7'h0 : _GEN_2931; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2933 = 10'h275 == io_inputs_1 ? 7'h0 : _GEN_2932; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2934 = 10'h276 == io_inputs_1 ? 7'h0 : _GEN_2933; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2935 = 10'h277 == io_inputs_1 ? 7'h0 : _GEN_2934; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2936 = 10'h278 == io_inputs_1 ? 7'h0 : _GEN_2935; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2937 = 10'h279 == io_inputs_1 ? 7'h0 : _GEN_2936; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2938 = 10'h27a == io_inputs_1 ? 7'h0 : _GEN_2937; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2939 = 10'h27b == io_inputs_1 ? 7'h0 : _GEN_2938; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2940 = 10'h27c == io_inputs_1 ? 7'h0 : _GEN_2939; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2941 = 10'h27d == io_inputs_1 ? 7'h0 : _GEN_2940; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2942 = 10'h27e == io_inputs_1 ? 7'h0 : _GEN_2941; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2943 = 10'h27f == io_inputs_1 ? 7'h0 : _GEN_2942; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2944 = 10'h280 == io_inputs_1 ? 7'h0 : _GEN_2943; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2945 = 10'h281 == io_inputs_1 ? 7'h0 : _GEN_2944; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2946 = 10'h282 == io_inputs_1 ? 7'h0 : _GEN_2945; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2947 = 10'h283 == io_inputs_1 ? 7'h0 : _GEN_2946; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2948 = 10'h284 == io_inputs_1 ? 7'h0 : _GEN_2947; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2949 = 10'h285 == io_inputs_1 ? 7'h0 : _GEN_2948; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2950 = 10'h286 == io_inputs_1 ? 7'h0 : _GEN_2949; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2951 = 10'h287 == io_inputs_1 ? 7'h0 : _GEN_2950; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2952 = 10'h288 == io_inputs_1 ? 7'h0 : _GEN_2951; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2953 = 10'h289 == io_inputs_1 ? 7'h0 : _GEN_2952; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2954 = 10'h28a == io_inputs_1 ? 7'h0 : _GEN_2953; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2955 = 10'h28b == io_inputs_1 ? 7'h0 : _GEN_2954; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2956 = 10'h28c == io_inputs_1 ? 7'h0 : _GEN_2955; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2957 = 10'h28d == io_inputs_1 ? 7'h0 : _GEN_2956; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2958 = 10'h28e == io_inputs_1 ? 7'h0 : _GEN_2957; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2959 = 10'h28f == io_inputs_1 ? 7'h0 : _GEN_2958; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2960 = 10'h290 == io_inputs_1 ? 7'h0 : _GEN_2959; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2961 = 10'h291 == io_inputs_1 ? 7'h0 : _GEN_2960; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2962 = 10'h292 == io_inputs_1 ? 7'h0 : _GEN_2961; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2963 = 10'h293 == io_inputs_1 ? 7'h0 : _GEN_2962; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2964 = 10'h294 == io_inputs_1 ? 7'h0 : _GEN_2963; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2965 = 10'h295 == io_inputs_1 ? 7'h0 : _GEN_2964; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2966 = 10'h296 == io_inputs_1 ? 7'h0 : _GEN_2965; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2967 = 10'h297 == io_inputs_1 ? 7'h0 : _GEN_2966; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2968 = 10'h298 == io_inputs_1 ? 7'h0 : _GEN_2967; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2969 = 10'h299 == io_inputs_1 ? 7'h0 : _GEN_2968; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2970 = 10'h29a == io_inputs_1 ? 7'h0 : _GEN_2969; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2971 = 10'h29b == io_inputs_1 ? 7'h0 : _GEN_2970; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2972 = 10'h29c == io_inputs_1 ? 7'h0 : _GEN_2971; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2973 = 10'h29d == io_inputs_1 ? 7'h0 : _GEN_2972; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2974 = 10'h29e == io_inputs_1 ? 7'h0 : _GEN_2973; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2975 = 10'h29f == io_inputs_1 ? 7'h0 : _GEN_2974; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2976 = 10'h2a0 == io_inputs_1 ? 7'h0 : _GEN_2975; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2977 = 10'h2a1 == io_inputs_1 ? 7'h0 : _GEN_2976; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2978 = 10'h2a2 == io_inputs_1 ? 7'h0 : _GEN_2977; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2979 = 10'h2a3 == io_inputs_1 ? 7'h0 : _GEN_2978; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2980 = 10'h2a4 == io_inputs_1 ? 7'h0 : _GEN_2979; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2981 = 10'h2a5 == io_inputs_1 ? 7'h0 : _GEN_2980; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2982 = 10'h2a6 == io_inputs_1 ? 7'h0 : _GEN_2981; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2983 = 10'h2a7 == io_inputs_1 ? 7'h0 : _GEN_2982; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2984 = 10'h2a8 == io_inputs_1 ? 7'h0 : _GEN_2983; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2985 = 10'h2a9 == io_inputs_1 ? 7'h0 : _GEN_2984; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2986 = 10'h2aa == io_inputs_1 ? 7'h0 : _GEN_2985; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2987 = 10'h2ab == io_inputs_1 ? 7'h0 : _GEN_2986; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2988 = 10'h2ac == io_inputs_1 ? 7'h0 : _GEN_2987; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2989 = 10'h2ad == io_inputs_1 ? 7'h0 : _GEN_2988; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2990 = 10'h2ae == io_inputs_1 ? 7'h0 : _GEN_2989; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2991 = 10'h2af == io_inputs_1 ? 7'h0 : _GEN_2990; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2992 = 10'h2b0 == io_inputs_1 ? 7'h0 : _GEN_2991; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2993 = 10'h2b1 == io_inputs_1 ? 7'h0 : _GEN_2992; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2994 = 10'h2b2 == io_inputs_1 ? 7'h0 : _GEN_2993; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2995 = 10'h2b3 == io_inputs_1 ? 7'h0 : _GEN_2994; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2996 = 10'h2b4 == io_inputs_1 ? 7'h0 : _GEN_2995; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2997 = 10'h2b5 == io_inputs_1 ? 7'h0 : _GEN_2996; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2998 = 10'h2b6 == io_inputs_1 ? 7'h0 : _GEN_2997; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_2999 = 10'h2b7 == io_inputs_1 ? 7'h0 : _GEN_2998; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3000 = 10'h2b8 == io_inputs_1 ? 7'h0 : _GEN_2999; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3001 = 10'h2b9 == io_inputs_1 ? 7'h0 : _GEN_3000; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3002 = 10'h2ba == io_inputs_1 ? 7'h0 : _GEN_3001; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3003 = 10'h2bb == io_inputs_1 ? 7'h0 : _GEN_3002; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3004 = 10'h2bc == io_inputs_1 ? 7'h0 : _GEN_3003; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3005 = 10'h2bd == io_inputs_1 ? 7'h0 : _GEN_3004; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3006 = 10'h2be == io_inputs_1 ? 7'h0 : _GEN_3005; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3007 = 10'h2bf == io_inputs_1 ? 7'h0 : _GEN_3006; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3008 = 10'h2c0 == io_inputs_1 ? 7'h0 : _GEN_3007; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3009 = 10'h2c1 == io_inputs_1 ? 7'h0 : _GEN_3008; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3010 = 10'h2c2 == io_inputs_1 ? 7'h0 : _GEN_3009; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3011 = 10'h2c3 == io_inputs_1 ? 7'h0 : _GEN_3010; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3012 = 10'h2c4 == io_inputs_1 ? 7'h0 : _GEN_3011; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3013 = 10'h2c5 == io_inputs_1 ? 7'h0 : _GEN_3012; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3014 = 10'h2c6 == io_inputs_1 ? 7'h0 : _GEN_3013; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3015 = 10'h2c7 == io_inputs_1 ? 7'h0 : _GEN_3014; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3016 = 10'h2c8 == io_inputs_1 ? 7'h0 : _GEN_3015; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3017 = 10'h2c9 == io_inputs_1 ? 7'h0 : _GEN_3016; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3018 = 10'h2ca == io_inputs_1 ? 7'h0 : _GEN_3017; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3019 = 10'h2cb == io_inputs_1 ? 7'h0 : _GEN_3018; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3020 = 10'h2cc == io_inputs_1 ? 7'h0 : _GEN_3019; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3021 = 10'h2cd == io_inputs_1 ? 7'h0 : _GEN_3020; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3022 = 10'h2ce == io_inputs_1 ? 7'h0 : _GEN_3021; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3023 = 10'h2cf == io_inputs_1 ? 7'h0 : _GEN_3022; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3024 = 10'h2d0 == io_inputs_1 ? 7'h0 : _GEN_3023; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3025 = 10'h2d1 == io_inputs_1 ? 7'h0 : _GEN_3024; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3026 = 10'h2d2 == io_inputs_1 ? 7'h0 : _GEN_3025; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3027 = 10'h2d3 == io_inputs_1 ? 7'h0 : _GEN_3026; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3028 = 10'h2d4 == io_inputs_1 ? 7'h0 : _GEN_3027; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3029 = 10'h2d5 == io_inputs_1 ? 7'h0 : _GEN_3028; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3030 = 10'h2d6 == io_inputs_1 ? 7'h0 : _GEN_3029; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3031 = 10'h2d7 == io_inputs_1 ? 7'h0 : _GEN_3030; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3032 = 10'h2d8 == io_inputs_1 ? 7'h0 : _GEN_3031; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3033 = 10'h2d9 == io_inputs_1 ? 7'h0 : _GEN_3032; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3034 = 10'h2da == io_inputs_1 ? 7'h0 : _GEN_3033; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3035 = 10'h2db == io_inputs_1 ? 7'h0 : _GEN_3034; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3036 = 10'h2dc == io_inputs_1 ? 7'h0 : _GEN_3035; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3037 = 10'h2dd == io_inputs_1 ? 7'h0 : _GEN_3036; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3038 = 10'h2de == io_inputs_1 ? 7'h0 : _GEN_3037; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3039 = 10'h2df == io_inputs_1 ? 7'h0 : _GEN_3038; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3040 = 10'h2e0 == io_inputs_1 ? 7'h0 : _GEN_3039; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3041 = 10'h2e1 == io_inputs_1 ? 7'h0 : _GEN_3040; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3042 = 10'h2e2 == io_inputs_1 ? 7'h0 : _GEN_3041; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3043 = 10'h2e3 == io_inputs_1 ? 7'h0 : _GEN_3042; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3044 = 10'h2e4 == io_inputs_1 ? 7'h0 : _GEN_3043; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3045 = 10'h2e5 == io_inputs_1 ? 7'h0 : _GEN_3044; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3046 = 10'h2e6 == io_inputs_1 ? 7'h0 : _GEN_3045; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3047 = 10'h2e7 == io_inputs_1 ? 7'h0 : _GEN_3046; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3048 = 10'h2e8 == io_inputs_1 ? 7'h0 : _GEN_3047; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3049 = 10'h2e9 == io_inputs_1 ? 7'h0 : _GEN_3048; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3050 = 10'h2ea == io_inputs_1 ? 7'h0 : _GEN_3049; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3051 = 10'h2eb == io_inputs_1 ? 7'h0 : _GEN_3050; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3052 = 10'h2ec == io_inputs_1 ? 7'h0 : _GEN_3051; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3053 = 10'h2ed == io_inputs_1 ? 7'h0 : _GEN_3052; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3054 = 10'h2ee == io_inputs_1 ? 7'h0 : _GEN_3053; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3055 = 10'h2ef == io_inputs_1 ? 7'h0 : _GEN_3054; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3056 = 10'h2f0 == io_inputs_1 ? 7'h0 : _GEN_3055; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3057 = 10'h2f1 == io_inputs_1 ? 7'h0 : _GEN_3056; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3058 = 10'h2f2 == io_inputs_1 ? 7'h0 : _GEN_3057; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3059 = 10'h2f3 == io_inputs_1 ? 7'h0 : _GEN_3058; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3060 = 10'h2f4 == io_inputs_1 ? 7'h0 : _GEN_3059; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3061 = 10'h2f5 == io_inputs_1 ? 7'h0 : _GEN_3060; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3062 = 10'h2f6 == io_inputs_1 ? 7'h0 : _GEN_3061; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3063 = 10'h2f7 == io_inputs_1 ? 7'h0 : _GEN_3062; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3064 = 10'h2f8 == io_inputs_1 ? 7'h0 : _GEN_3063; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3065 = 10'h2f9 == io_inputs_1 ? 7'h0 : _GEN_3064; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3066 = 10'h2fa == io_inputs_1 ? 7'h0 : _GEN_3065; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3067 = 10'h2fb == io_inputs_1 ? 7'h0 : _GEN_3066; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3068 = 10'h2fc == io_inputs_1 ? 7'h0 : _GEN_3067; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3069 = 10'h2fd == io_inputs_1 ? 7'h0 : _GEN_3068; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3070 = 10'h2fe == io_inputs_1 ? 7'h0 : _GEN_3069; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3071 = 10'h2ff == io_inputs_1 ? 7'h0 : _GEN_3070; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3072 = 10'h300 == io_inputs_1 ? 7'h0 : _GEN_3071; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3073 = 10'h301 == io_inputs_1 ? 7'h0 : _GEN_3072; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3074 = 10'h302 == io_inputs_1 ? 7'h0 : _GEN_3073; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3075 = 10'h303 == io_inputs_1 ? 7'h0 : _GEN_3074; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3076 = 10'h304 == io_inputs_1 ? 7'h0 : _GEN_3075; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3077 = 10'h305 == io_inputs_1 ? 7'h0 : _GEN_3076; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3078 = 10'h306 == io_inputs_1 ? 7'h0 : _GEN_3077; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3079 = 10'h307 == io_inputs_1 ? 7'h0 : _GEN_3078; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3080 = 10'h308 == io_inputs_1 ? 7'h0 : _GEN_3079; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3081 = 10'h309 == io_inputs_1 ? 7'h0 : _GEN_3080; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3082 = 10'h30a == io_inputs_1 ? 7'h0 : _GEN_3081; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3083 = 10'h30b == io_inputs_1 ? 7'h0 : _GEN_3082; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3084 = 10'h30c == io_inputs_1 ? 7'h0 : _GEN_3083; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3085 = 10'h30d == io_inputs_1 ? 7'h0 : _GEN_3084; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3086 = 10'h30e == io_inputs_1 ? 7'h0 : _GEN_3085; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3087 = 10'h30f == io_inputs_1 ? 7'h0 : _GEN_3086; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3088 = 10'h310 == io_inputs_1 ? 7'h0 : _GEN_3087; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3089 = 10'h311 == io_inputs_1 ? 7'h0 : _GEN_3088; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3090 = 10'h312 == io_inputs_1 ? 7'h0 : _GEN_3089; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3091 = 10'h313 == io_inputs_1 ? 7'h0 : _GEN_3090; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3092 = 10'h314 == io_inputs_1 ? 7'h0 : _GEN_3091; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3093 = 10'h315 == io_inputs_1 ? 7'h0 : _GEN_3092; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3094 = 10'h316 == io_inputs_1 ? 7'h0 : _GEN_3093; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3095 = 10'h317 == io_inputs_1 ? 7'h0 : _GEN_3094; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3096 = 10'h318 == io_inputs_1 ? 7'h0 : _GEN_3095; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3097 = 10'h319 == io_inputs_1 ? 7'h0 : _GEN_3096; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3098 = 10'h31a == io_inputs_1 ? 7'h0 : _GEN_3097; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3099 = 10'h31b == io_inputs_1 ? 7'h0 : _GEN_3098; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3100 = 10'h31c == io_inputs_1 ? 7'h0 : _GEN_3099; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3101 = 10'h31d == io_inputs_1 ? 7'h0 : _GEN_3100; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3102 = 10'h31e == io_inputs_1 ? 7'h0 : _GEN_3101; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3103 = 10'h31f == io_inputs_1 ? 7'h0 : _GEN_3102; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3104 = 10'h320 == io_inputs_1 ? 7'h0 : _GEN_3103; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3105 = 10'h321 == io_inputs_1 ? 7'h0 : _GEN_3104; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3106 = 10'h322 == io_inputs_1 ? 7'h0 : _GEN_3105; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3107 = 10'h323 == io_inputs_1 ? 7'h0 : _GEN_3106; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3108 = 10'h324 == io_inputs_1 ? 7'h0 : _GEN_3107; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3109 = 10'h325 == io_inputs_1 ? 7'h0 : _GEN_3108; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3110 = 10'h326 == io_inputs_1 ? 7'h0 : _GEN_3109; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3111 = 10'h327 == io_inputs_1 ? 7'h0 : _GEN_3110; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3112 = 10'h328 == io_inputs_1 ? 7'h0 : _GEN_3111; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3113 = 10'h329 == io_inputs_1 ? 7'h0 : _GEN_3112; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3114 = 10'h32a == io_inputs_1 ? 7'h0 : _GEN_3113; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3115 = 10'h32b == io_inputs_1 ? 7'h0 : _GEN_3114; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3116 = 10'h32c == io_inputs_1 ? 7'h0 : _GEN_3115; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3117 = 10'h32d == io_inputs_1 ? 7'h0 : _GEN_3116; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3118 = 10'h32e == io_inputs_1 ? 7'h0 : _GEN_3117; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3119 = 10'h32f == io_inputs_1 ? 7'h0 : _GEN_3118; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3120 = 10'h330 == io_inputs_1 ? 7'h0 : _GEN_3119; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3121 = 10'h331 == io_inputs_1 ? 7'h0 : _GEN_3120; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3122 = 10'h332 == io_inputs_1 ? 7'h0 : _GEN_3121; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3123 = 10'h333 == io_inputs_1 ? 7'h0 : _GEN_3122; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3124 = 10'h334 == io_inputs_1 ? 7'h0 : _GEN_3123; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3125 = 10'h335 == io_inputs_1 ? 7'h0 : _GEN_3124; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3126 = 10'h336 == io_inputs_1 ? 7'h0 : _GEN_3125; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3127 = 10'h337 == io_inputs_1 ? 7'h0 : _GEN_3126; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3128 = 10'h338 == io_inputs_1 ? 7'h0 : _GEN_3127; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3129 = 10'h339 == io_inputs_1 ? 7'h0 : _GEN_3128; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3130 = 10'h33a == io_inputs_1 ? 7'h0 : _GEN_3129; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3131 = 10'h33b == io_inputs_1 ? 7'h0 : _GEN_3130; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3132 = 10'h33c == io_inputs_1 ? 7'h0 : _GEN_3131; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3133 = 10'h33d == io_inputs_1 ? 7'h0 : _GEN_3132; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3134 = 10'h33e == io_inputs_1 ? 7'h0 : _GEN_3133; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3135 = 10'h33f == io_inputs_1 ? 7'h0 : _GEN_3134; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3136 = 10'h340 == io_inputs_1 ? 7'h0 : _GEN_3135; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3137 = 10'h341 == io_inputs_1 ? 7'h0 : _GEN_3136; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3138 = 10'h342 == io_inputs_1 ? 7'h0 : _GEN_3137; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3139 = 10'h343 == io_inputs_1 ? 7'h0 : _GEN_3138; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3140 = 10'h344 == io_inputs_1 ? 7'h0 : _GEN_3139; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3141 = 10'h345 == io_inputs_1 ? 7'h0 : _GEN_3140; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3142 = 10'h346 == io_inputs_1 ? 7'h0 : _GEN_3141; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3143 = 10'h347 == io_inputs_1 ? 7'h0 : _GEN_3142; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3144 = 10'h348 == io_inputs_1 ? 7'h0 : _GEN_3143; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3145 = 10'h349 == io_inputs_1 ? 7'h0 : _GEN_3144; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3146 = 10'h34a == io_inputs_1 ? 7'h0 : _GEN_3145; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3147 = 10'h34b == io_inputs_1 ? 7'h0 : _GEN_3146; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3148 = 10'h34c == io_inputs_1 ? 7'h0 : _GEN_3147; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3149 = 10'h34d == io_inputs_1 ? 7'h0 : _GEN_3148; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3150 = 10'h34e == io_inputs_1 ? 7'h0 : _GEN_3149; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3151 = 10'h34f == io_inputs_1 ? 7'h0 : _GEN_3150; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3152 = 10'h350 == io_inputs_1 ? 7'h0 : _GEN_3151; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3153 = 10'h351 == io_inputs_1 ? 7'h0 : _GEN_3152; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3154 = 10'h352 == io_inputs_1 ? 7'h0 : _GEN_3153; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3155 = 10'h353 == io_inputs_1 ? 7'h0 : _GEN_3154; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3156 = 10'h354 == io_inputs_1 ? 7'h0 : _GEN_3155; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3157 = 10'h355 == io_inputs_1 ? 7'h0 : _GEN_3156; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3158 = 10'h356 == io_inputs_1 ? 7'h0 : _GEN_3157; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3159 = 10'h357 == io_inputs_1 ? 7'h0 : _GEN_3158; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3160 = 10'h358 == io_inputs_1 ? 7'h0 : _GEN_3159; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3161 = 10'h359 == io_inputs_1 ? 7'h0 : _GEN_3160; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3162 = 10'h35a == io_inputs_1 ? 7'h0 : _GEN_3161; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3163 = 10'h35b == io_inputs_1 ? 7'h0 : _GEN_3162; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3164 = 10'h35c == io_inputs_1 ? 7'h0 : _GEN_3163; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3165 = 10'h35d == io_inputs_1 ? 7'h0 : _GEN_3164; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3166 = 10'h35e == io_inputs_1 ? 7'h0 : _GEN_3165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3167 = 10'h35f == io_inputs_1 ? 7'h0 : _GEN_3166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3168 = 10'h360 == io_inputs_1 ? 7'h0 : _GEN_3167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3169 = 10'h361 == io_inputs_1 ? 7'h0 : _GEN_3168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3170 = 10'h362 == io_inputs_1 ? 7'h0 : _GEN_3169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3171 = 10'h363 == io_inputs_1 ? 7'h0 : _GEN_3170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3172 = 10'h364 == io_inputs_1 ? 7'h0 : _GEN_3171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3173 = 10'h365 == io_inputs_1 ? 7'h0 : _GEN_3172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3174 = 10'h366 == io_inputs_1 ? 7'h0 : _GEN_3173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3175 = 10'h367 == io_inputs_1 ? 7'h0 : _GEN_3174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3176 = 10'h368 == io_inputs_1 ? 7'h0 : _GEN_3175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3177 = 10'h369 == io_inputs_1 ? 7'h0 : _GEN_3176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3178 = 10'h36a == io_inputs_1 ? 7'h0 : _GEN_3177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3179 = 10'h36b == io_inputs_1 ? 7'h0 : _GEN_3178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3180 = 10'h36c == io_inputs_1 ? 7'h0 : _GEN_3179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3181 = 10'h36d == io_inputs_1 ? 7'h0 : _GEN_3180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3182 = 10'h36e == io_inputs_1 ? 7'h0 : _GEN_3181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3183 = 10'h36f == io_inputs_1 ? 7'h0 : _GEN_3182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3184 = 10'h370 == io_inputs_1 ? 7'h0 : _GEN_3183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3185 = 10'h371 == io_inputs_1 ? 7'h0 : _GEN_3184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3186 = 10'h372 == io_inputs_1 ? 7'h0 : _GEN_3185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3187 = 10'h373 == io_inputs_1 ? 7'h0 : _GEN_3186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3188 = 10'h374 == io_inputs_1 ? 7'h0 : _GEN_3187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3189 = 10'h375 == io_inputs_1 ? 7'h0 : _GEN_3188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3190 = 10'h376 == io_inputs_1 ? 7'h0 : _GEN_3189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3191 = 10'h377 == io_inputs_1 ? 7'h0 : _GEN_3190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3192 = 10'h378 == io_inputs_1 ? 7'h0 : _GEN_3191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3193 = 10'h379 == io_inputs_1 ? 7'h0 : _GEN_3192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3194 = 10'h37a == io_inputs_1 ? 7'h0 : _GEN_3193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3195 = 10'h37b == io_inputs_1 ? 7'h0 : _GEN_3194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3196 = 10'h37c == io_inputs_1 ? 7'h0 : _GEN_3195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3197 = 10'h37d == io_inputs_1 ? 7'h0 : _GEN_3196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3198 = 10'h37e == io_inputs_1 ? 7'h0 : _GEN_3197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3199 = 10'h37f == io_inputs_1 ? 7'h0 : _GEN_3198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3200 = 10'h380 == io_inputs_1 ? 7'h0 : _GEN_3199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3201 = 10'h381 == io_inputs_1 ? 7'h0 : _GEN_3200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3202 = 10'h382 == io_inputs_1 ? 7'h0 : _GEN_3201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3203 = 10'h383 == io_inputs_1 ? 7'h0 : _GEN_3202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3204 = 10'h384 == io_inputs_1 ? 7'h0 : _GEN_3203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3205 = 10'h385 == io_inputs_1 ? 7'h0 : _GEN_3204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3206 = 10'h386 == io_inputs_1 ? 7'h0 : _GEN_3205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3207 = 10'h387 == io_inputs_1 ? 7'h0 : _GEN_3206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3208 = 10'h388 == io_inputs_1 ? 7'h0 : _GEN_3207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3209 = 10'h389 == io_inputs_1 ? 7'h0 : _GEN_3208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3210 = 10'h38a == io_inputs_1 ? 7'h0 : _GEN_3209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3211 = 10'h38b == io_inputs_1 ? 7'h0 : _GEN_3210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3212 = 10'h38c == io_inputs_1 ? 7'h0 : _GEN_3211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3213 = 10'h38d == io_inputs_1 ? 7'h0 : _GEN_3212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3214 = 10'h38e == io_inputs_1 ? 7'h0 : _GEN_3213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3215 = 10'h38f == io_inputs_1 ? 7'h0 : _GEN_3214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3216 = 10'h390 == io_inputs_1 ? 7'h0 : _GEN_3215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3217 = 10'h391 == io_inputs_1 ? 7'h0 : _GEN_3216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3218 = 10'h392 == io_inputs_1 ? 7'h0 : _GEN_3217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3219 = 10'h393 == io_inputs_1 ? 7'h0 : _GEN_3218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3220 = 10'h394 == io_inputs_1 ? 7'h0 : _GEN_3219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3221 = 10'h395 == io_inputs_1 ? 7'h0 : _GEN_3220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3222 = 10'h396 == io_inputs_1 ? 7'h0 : _GEN_3221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3223 = 10'h397 == io_inputs_1 ? 7'h0 : _GEN_3222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3224 = 10'h398 == io_inputs_1 ? 7'h0 : _GEN_3223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3225 = 10'h399 == io_inputs_1 ? 7'h0 : _GEN_3224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3226 = 10'h39a == io_inputs_1 ? 7'h0 : _GEN_3225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3227 = 10'h39b == io_inputs_1 ? 7'h0 : _GEN_3226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3228 = 10'h39c == io_inputs_1 ? 7'h0 : _GEN_3227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3229 = 10'h39d == io_inputs_1 ? 7'h0 : _GEN_3228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3230 = 10'h39e == io_inputs_1 ? 7'h0 : _GEN_3229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3231 = 10'h39f == io_inputs_1 ? 7'h0 : _GEN_3230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3232 = 10'h3a0 == io_inputs_1 ? 7'h0 : _GEN_3231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3233 = 10'h3a1 == io_inputs_1 ? 7'h0 : _GEN_3232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3234 = 10'h3a2 == io_inputs_1 ? 7'h0 : _GEN_3233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3235 = 10'h3a3 == io_inputs_1 ? 7'h0 : _GEN_3234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3236 = 10'h3a4 == io_inputs_1 ? 7'h0 : _GEN_3235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3237 = 10'h3a5 == io_inputs_1 ? 7'h0 : _GEN_3236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3238 = 10'h3a6 == io_inputs_1 ? 7'h0 : _GEN_3237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3239 = 10'h3a7 == io_inputs_1 ? 7'h0 : _GEN_3238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3240 = 10'h3a8 == io_inputs_1 ? 7'h0 : _GEN_3239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3241 = 10'h3a9 == io_inputs_1 ? 7'h0 : _GEN_3240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3242 = 10'h3aa == io_inputs_1 ? 7'h0 : _GEN_3241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3243 = 10'h3ab == io_inputs_1 ? 7'h0 : _GEN_3242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3244 = 10'h3ac == io_inputs_1 ? 7'h0 : _GEN_3243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3245 = 10'h3ad == io_inputs_1 ? 7'h0 : _GEN_3244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3246 = 10'h3ae == io_inputs_1 ? 7'h0 : _GEN_3245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3247 = 10'h3af == io_inputs_1 ? 7'h0 : _GEN_3246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3248 = 10'h3b0 == io_inputs_1 ? 7'h0 : _GEN_3247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3249 = 10'h3b1 == io_inputs_1 ? 7'h0 : _GEN_3248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3250 = 10'h3b2 == io_inputs_1 ? 7'h0 : _GEN_3249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3251 = 10'h3b3 == io_inputs_1 ? 7'h0 : _GEN_3250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3252 = 10'h3b4 == io_inputs_1 ? 7'h0 : _GEN_3251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3253 = 10'h3b5 == io_inputs_1 ? 7'h0 : _GEN_3252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3254 = 10'h3b6 == io_inputs_1 ? 7'h0 : _GEN_3253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3255 = 10'h3b7 == io_inputs_1 ? 7'h0 : _GEN_3254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3256 = 10'h3b8 == io_inputs_1 ? 7'h0 : _GEN_3255; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3257 = 10'h3b9 == io_inputs_1 ? 7'h0 : _GEN_3256; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3258 = 10'h3ba == io_inputs_1 ? 7'h0 : _GEN_3257; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3259 = 10'h3bb == io_inputs_1 ? 7'h0 : _GEN_3258; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3260 = 10'h3bc == io_inputs_1 ? 7'h0 : _GEN_3259; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3261 = 10'h3bd == io_inputs_1 ? 7'h0 : _GEN_3260; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3262 = 10'h3be == io_inputs_1 ? 7'h0 : _GEN_3261; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3263 = 10'h3bf == io_inputs_1 ? 7'h0 : _GEN_3262; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3264 = 10'h3c0 == io_inputs_1 ? 7'h0 : _GEN_3263; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3265 = 10'h3c1 == io_inputs_1 ? 7'h0 : _GEN_3264; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3266 = 10'h3c2 == io_inputs_1 ? 7'h0 : _GEN_3265; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3267 = 10'h3c3 == io_inputs_1 ? 7'h0 : _GEN_3266; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3268 = 10'h3c4 == io_inputs_1 ? 7'h0 : _GEN_3267; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3269 = 10'h3c5 == io_inputs_1 ? 7'h0 : _GEN_3268; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3270 = 10'h3c6 == io_inputs_1 ? 7'h0 : _GEN_3269; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3271 = 10'h3c7 == io_inputs_1 ? 7'h0 : _GEN_3270; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3272 = 10'h3c8 == io_inputs_1 ? 7'h0 : _GEN_3271; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3273 = 10'h3c9 == io_inputs_1 ? 7'h0 : _GEN_3272; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3274 = 10'h3ca == io_inputs_1 ? 7'h0 : _GEN_3273; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3275 = 10'h3cb == io_inputs_1 ? 7'h0 : _GEN_3274; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3276 = 10'h3cc == io_inputs_1 ? 7'h0 : _GEN_3275; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3277 = 10'h3cd == io_inputs_1 ? 7'h0 : _GEN_3276; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3278 = 10'h3ce == io_inputs_1 ? 7'h0 : _GEN_3277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3279 = 10'h3cf == io_inputs_1 ? 7'h0 : _GEN_3278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3280 = 10'h3d0 == io_inputs_1 ? 7'h0 : _GEN_3279; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3281 = 10'h3d1 == io_inputs_1 ? 7'h0 : _GEN_3280; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3282 = 10'h3d2 == io_inputs_1 ? 7'h0 : _GEN_3281; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3283 = 10'h3d3 == io_inputs_1 ? 7'h0 : _GEN_3282; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3284 = 10'h3d4 == io_inputs_1 ? 7'h0 : _GEN_3283; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3285 = 10'h3d5 == io_inputs_1 ? 7'h0 : _GEN_3284; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3286 = 10'h3d6 == io_inputs_1 ? 7'h0 : _GEN_3285; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3287 = 10'h3d7 == io_inputs_1 ? 7'h0 : _GEN_3286; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3288 = 10'h3d8 == io_inputs_1 ? 7'h0 : _GEN_3287; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3289 = 10'h3d9 == io_inputs_1 ? 7'h0 : _GEN_3288; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3290 = 10'h3da == io_inputs_1 ? 7'h0 : _GEN_3289; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3291 = 10'h3db == io_inputs_1 ? 7'h0 : _GEN_3290; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3292 = 10'h3dc == io_inputs_1 ? 7'h0 : _GEN_3291; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3293 = 10'h3dd == io_inputs_1 ? 7'h0 : _GEN_3292; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3294 = 10'h3de == io_inputs_1 ? 7'h0 : _GEN_3293; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3295 = 10'h3df == io_inputs_1 ? 7'h0 : _GEN_3294; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3296 = 10'h3e0 == io_inputs_1 ? 7'h0 : _GEN_3295; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3297 = 10'h3e1 == io_inputs_1 ? 7'h0 : _GEN_3296; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3298 = 10'h3e2 == io_inputs_1 ? 7'h0 : _GEN_3297; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3299 = 10'h3e3 == io_inputs_1 ? 7'h0 : _GEN_3298; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3300 = 10'h3e4 == io_inputs_1 ? 7'h0 : _GEN_3299; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3301 = 10'h3e5 == io_inputs_1 ? 7'h0 : _GEN_3300; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3302 = 10'h3e6 == io_inputs_1 ? 7'h0 : _GEN_3301; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3303 = 10'h3e7 == io_inputs_1 ? 7'h0 : _GEN_3302; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3304 = 10'h3e8 == io_inputs_1 ? 7'h0 : _GEN_3303; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3305 = 10'h3e9 == io_inputs_1 ? 7'h0 : _GEN_3304; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3306 = 10'h3ea == io_inputs_1 ? 7'h0 : _GEN_3305; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3307 = 10'h3eb == io_inputs_1 ? 7'h0 : _GEN_3306; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3308 = 10'h3ec == io_inputs_1 ? 7'h0 : _GEN_3307; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3309 = 10'h3ed == io_inputs_1 ? 7'h0 : _GEN_3308; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3310 = 10'h3ee == io_inputs_1 ? 7'h0 : _GEN_3309; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3311 = 10'h3ef == io_inputs_1 ? 7'h0 : _GEN_3310; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3312 = 10'h3f0 == io_inputs_1 ? 7'h0 : _GEN_3311; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3313 = 10'h3f1 == io_inputs_1 ? 7'h0 : _GEN_3312; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3314 = 10'h3f2 == io_inputs_1 ? 7'h0 : _GEN_3313; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3315 = 10'h3f3 == io_inputs_1 ? 7'h0 : _GEN_3314; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3316 = 10'h3f4 == io_inputs_1 ? 7'h0 : _GEN_3315; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3317 = 10'h3f5 == io_inputs_1 ? 7'h0 : _GEN_3316; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3318 = 10'h3f6 == io_inputs_1 ? 7'h0 : _GEN_3317; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3319 = 10'h3f7 == io_inputs_1 ? 7'h0 : _GEN_3318; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3320 = 10'h3f8 == io_inputs_1 ? 7'h0 : _GEN_3319; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3321 = 10'h3f9 == io_inputs_1 ? 7'h0 : _GEN_3320; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3322 = 10'h3fa == io_inputs_1 ? 7'h0 : _GEN_3321; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3323 = 10'h3fb == io_inputs_1 ? 7'h0 : _GEN_3322; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3324 = 10'h3fc == io_inputs_1 ? 7'h0 : _GEN_3323; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3325 = 10'h3fd == io_inputs_1 ? 7'h0 : _GEN_3324; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3326 = 10'h3fe == io_inputs_1 ? 7'h0 : _GEN_3325; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3327 = 10'h3ff == io_inputs_1 ? 7'h0 : _GEN_3326; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3529 = 10'hc9 == io_inputs_1 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3530 = 10'hca == io_inputs_1 ? 7'h2 : _GEN_3529; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3531 = 10'hcb == io_inputs_1 ? 7'h3 : _GEN_3530; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3532 = 10'hcc == io_inputs_1 ? 7'h4 : _GEN_3531; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3533 = 10'hcd == io_inputs_1 ? 7'h5 : _GEN_3532; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3534 = 10'hce == io_inputs_1 ? 7'h6 : _GEN_3533; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3535 = 10'hcf == io_inputs_1 ? 7'h7 : _GEN_3534; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3536 = 10'hd0 == io_inputs_1 ? 7'h8 : _GEN_3535; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3537 = 10'hd1 == io_inputs_1 ? 7'h9 : _GEN_3536; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3538 = 10'hd2 == io_inputs_1 ? 7'ha : _GEN_3537; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3539 = 10'hd3 == io_inputs_1 ? 7'hb : _GEN_3538; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3540 = 10'hd4 == io_inputs_1 ? 7'hc : _GEN_3539; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3541 = 10'hd5 == io_inputs_1 ? 7'hd : _GEN_3540; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3542 = 10'hd6 == io_inputs_1 ? 7'he : _GEN_3541; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3543 = 10'hd7 == io_inputs_1 ? 7'hf : _GEN_3542; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3544 = 10'hd8 == io_inputs_1 ? 7'h10 : _GEN_3543; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3545 = 10'hd9 == io_inputs_1 ? 7'h11 : _GEN_3544; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3546 = 10'hda == io_inputs_1 ? 7'h12 : _GEN_3545; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3547 = 10'hdb == io_inputs_1 ? 7'h13 : _GEN_3546; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3548 = 10'hdc == io_inputs_1 ? 7'h14 : _GEN_3547; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3549 = 10'hdd == io_inputs_1 ? 7'h15 : _GEN_3548; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3550 = 10'hde == io_inputs_1 ? 7'h16 : _GEN_3549; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3551 = 10'hdf == io_inputs_1 ? 7'h17 : _GEN_3550; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3552 = 10'he0 == io_inputs_1 ? 7'h18 : _GEN_3551; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3553 = 10'he1 == io_inputs_1 ? 7'h19 : _GEN_3552; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3554 = 10'he2 == io_inputs_1 ? 7'h1a : _GEN_3553; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3555 = 10'he3 == io_inputs_1 ? 7'h1b : _GEN_3554; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3556 = 10'he4 == io_inputs_1 ? 7'h1c : _GEN_3555; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3557 = 10'he5 == io_inputs_1 ? 7'h1d : _GEN_3556; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3558 = 10'he6 == io_inputs_1 ? 7'h1e : _GEN_3557; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3559 = 10'he7 == io_inputs_1 ? 7'h1f : _GEN_3558; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3560 = 10'he8 == io_inputs_1 ? 7'h20 : _GEN_3559; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3561 = 10'he9 == io_inputs_1 ? 7'h21 : _GEN_3560; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3562 = 10'hea == io_inputs_1 ? 7'h22 : _GEN_3561; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3563 = 10'heb == io_inputs_1 ? 7'h23 : _GEN_3562; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3564 = 10'hec == io_inputs_1 ? 7'h24 : _GEN_3563; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3565 = 10'hed == io_inputs_1 ? 7'h25 : _GEN_3564; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3566 = 10'hee == io_inputs_1 ? 7'h26 : _GEN_3565; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3567 = 10'hef == io_inputs_1 ? 7'h27 : _GEN_3566; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3568 = 10'hf0 == io_inputs_1 ? 7'h28 : _GEN_3567; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3569 = 10'hf1 == io_inputs_1 ? 7'h29 : _GEN_3568; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3570 = 10'hf2 == io_inputs_1 ? 7'h2a : _GEN_3569; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3571 = 10'hf3 == io_inputs_1 ? 7'h2b : _GEN_3570; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3572 = 10'hf4 == io_inputs_1 ? 7'h2c : _GEN_3571; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3573 = 10'hf5 == io_inputs_1 ? 7'h2d : _GEN_3572; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3574 = 10'hf6 == io_inputs_1 ? 7'h2e : _GEN_3573; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3575 = 10'hf7 == io_inputs_1 ? 7'h2f : _GEN_3574; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3576 = 10'hf8 == io_inputs_1 ? 7'h30 : _GEN_3575; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3577 = 10'hf9 == io_inputs_1 ? 7'h31 : _GEN_3576; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3578 = 10'hfa == io_inputs_1 ? 7'h32 : _GEN_3577; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3579 = 10'hfb == io_inputs_1 ? 7'h33 : _GEN_3578; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3580 = 10'hfc == io_inputs_1 ? 7'h34 : _GEN_3579; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3581 = 10'hfd == io_inputs_1 ? 7'h35 : _GEN_3580; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3582 = 10'hfe == io_inputs_1 ? 7'h36 : _GEN_3581; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3583 = 10'hff == io_inputs_1 ? 7'h37 : _GEN_3582; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3584 = 10'h100 == io_inputs_1 ? 7'h38 : _GEN_3583; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3585 = 10'h101 == io_inputs_1 ? 7'h39 : _GEN_3584; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3586 = 10'h102 == io_inputs_1 ? 7'h3a : _GEN_3585; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3587 = 10'h103 == io_inputs_1 ? 7'h3b : _GEN_3586; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3588 = 10'h104 == io_inputs_1 ? 7'h3c : _GEN_3587; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3589 = 10'h105 == io_inputs_1 ? 7'h3d : _GEN_3588; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3590 = 10'h106 == io_inputs_1 ? 7'h3e : _GEN_3589; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3591 = 10'h107 == io_inputs_1 ? 7'h3f : _GEN_3590; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3592 = 10'h108 == io_inputs_1 ? 7'h40 : _GEN_3591; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3593 = 10'h109 == io_inputs_1 ? 7'h41 : _GEN_3592; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3594 = 10'h10a == io_inputs_1 ? 7'h42 : _GEN_3593; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3595 = 10'h10b == io_inputs_1 ? 7'h43 : _GEN_3594; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3596 = 10'h10c == io_inputs_1 ? 7'h44 : _GEN_3595; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3597 = 10'h10d == io_inputs_1 ? 7'h45 : _GEN_3596; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3598 = 10'h10e == io_inputs_1 ? 7'h46 : _GEN_3597; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3599 = 10'h10f == io_inputs_1 ? 7'h47 : _GEN_3598; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3600 = 10'h110 == io_inputs_1 ? 7'h48 : _GEN_3599; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3601 = 10'h111 == io_inputs_1 ? 7'h49 : _GEN_3600; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3602 = 10'h112 == io_inputs_1 ? 7'h4a : _GEN_3601; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3603 = 10'h113 == io_inputs_1 ? 7'h4b : _GEN_3602; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3604 = 10'h114 == io_inputs_1 ? 7'h4c : _GEN_3603; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3605 = 10'h115 == io_inputs_1 ? 7'h4d : _GEN_3604; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3606 = 10'h116 == io_inputs_1 ? 7'h4e : _GEN_3605; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3607 = 10'h117 == io_inputs_1 ? 7'h4f : _GEN_3606; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3608 = 10'h118 == io_inputs_1 ? 7'h50 : _GEN_3607; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3609 = 10'h119 == io_inputs_1 ? 7'h51 : _GEN_3608; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3610 = 10'h11a == io_inputs_1 ? 7'h52 : _GEN_3609; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3611 = 10'h11b == io_inputs_1 ? 7'h53 : _GEN_3610; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3612 = 10'h11c == io_inputs_1 ? 7'h54 : _GEN_3611; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3613 = 10'h11d == io_inputs_1 ? 7'h55 : _GEN_3612; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3614 = 10'h11e == io_inputs_1 ? 7'h56 : _GEN_3613; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3615 = 10'h11f == io_inputs_1 ? 7'h57 : _GEN_3614; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3616 = 10'h120 == io_inputs_1 ? 7'h58 : _GEN_3615; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3617 = 10'h121 == io_inputs_1 ? 7'h59 : _GEN_3616; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3618 = 10'h122 == io_inputs_1 ? 7'h5a : _GEN_3617; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3619 = 10'h123 == io_inputs_1 ? 7'h5b : _GEN_3618; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3620 = 10'h124 == io_inputs_1 ? 7'h5c : _GEN_3619; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3621 = 10'h125 == io_inputs_1 ? 7'h5d : _GEN_3620; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3622 = 10'h126 == io_inputs_1 ? 7'h5e : _GEN_3621; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3623 = 10'h127 == io_inputs_1 ? 7'h5f : _GEN_3622; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3624 = 10'h128 == io_inputs_1 ? 7'h60 : _GEN_3623; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3625 = 10'h129 == io_inputs_1 ? 7'h61 : _GEN_3624; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3626 = 10'h12a == io_inputs_1 ? 7'h62 : _GEN_3625; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3627 = 10'h12b == io_inputs_1 ? 7'h63 : _GEN_3626; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3628 = 10'h12c == io_inputs_1 ? 7'h64 : _GEN_3627; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3629 = 10'h12d == io_inputs_1 ? 7'h0 : _GEN_3628; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3630 = 10'h12e == io_inputs_1 ? 7'h0 : _GEN_3629; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3631 = 10'h12f == io_inputs_1 ? 7'h0 : _GEN_3630; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3632 = 10'h130 == io_inputs_1 ? 7'h0 : _GEN_3631; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3633 = 10'h131 == io_inputs_1 ? 7'h0 : _GEN_3632; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3634 = 10'h132 == io_inputs_1 ? 7'h0 : _GEN_3633; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3635 = 10'h133 == io_inputs_1 ? 7'h0 : _GEN_3634; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3636 = 10'h134 == io_inputs_1 ? 7'h0 : _GEN_3635; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3637 = 10'h135 == io_inputs_1 ? 7'h0 : _GEN_3636; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3638 = 10'h136 == io_inputs_1 ? 7'h0 : _GEN_3637; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3639 = 10'h137 == io_inputs_1 ? 7'h0 : _GEN_3638; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3640 = 10'h138 == io_inputs_1 ? 7'h0 : _GEN_3639; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3641 = 10'h139 == io_inputs_1 ? 7'h0 : _GEN_3640; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3642 = 10'h13a == io_inputs_1 ? 7'h0 : _GEN_3641; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3643 = 10'h13b == io_inputs_1 ? 7'h0 : _GEN_3642; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3644 = 10'h13c == io_inputs_1 ? 7'h0 : _GEN_3643; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3645 = 10'h13d == io_inputs_1 ? 7'h0 : _GEN_3644; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3646 = 10'h13e == io_inputs_1 ? 7'h0 : _GEN_3645; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3647 = 10'h13f == io_inputs_1 ? 7'h0 : _GEN_3646; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3648 = 10'h140 == io_inputs_1 ? 7'h0 : _GEN_3647; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3649 = 10'h141 == io_inputs_1 ? 7'h0 : _GEN_3648; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3650 = 10'h142 == io_inputs_1 ? 7'h0 : _GEN_3649; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3651 = 10'h143 == io_inputs_1 ? 7'h0 : _GEN_3650; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3652 = 10'h144 == io_inputs_1 ? 7'h0 : _GEN_3651; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3653 = 10'h145 == io_inputs_1 ? 7'h0 : _GEN_3652; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3654 = 10'h146 == io_inputs_1 ? 7'h0 : _GEN_3653; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3655 = 10'h147 == io_inputs_1 ? 7'h0 : _GEN_3654; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3656 = 10'h148 == io_inputs_1 ? 7'h0 : _GEN_3655; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3657 = 10'h149 == io_inputs_1 ? 7'h0 : _GEN_3656; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3658 = 10'h14a == io_inputs_1 ? 7'h0 : _GEN_3657; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3659 = 10'h14b == io_inputs_1 ? 7'h0 : _GEN_3658; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3660 = 10'h14c == io_inputs_1 ? 7'h0 : _GEN_3659; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3661 = 10'h14d == io_inputs_1 ? 7'h0 : _GEN_3660; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3662 = 10'h14e == io_inputs_1 ? 7'h0 : _GEN_3661; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3663 = 10'h14f == io_inputs_1 ? 7'h0 : _GEN_3662; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3664 = 10'h150 == io_inputs_1 ? 7'h0 : _GEN_3663; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3665 = 10'h151 == io_inputs_1 ? 7'h0 : _GEN_3664; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3666 = 10'h152 == io_inputs_1 ? 7'h0 : _GEN_3665; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3667 = 10'h153 == io_inputs_1 ? 7'h0 : _GEN_3666; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3668 = 10'h154 == io_inputs_1 ? 7'h0 : _GEN_3667; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3669 = 10'h155 == io_inputs_1 ? 7'h0 : _GEN_3668; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3670 = 10'h156 == io_inputs_1 ? 7'h0 : _GEN_3669; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3671 = 10'h157 == io_inputs_1 ? 7'h0 : _GEN_3670; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3672 = 10'h158 == io_inputs_1 ? 7'h0 : _GEN_3671; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3673 = 10'h159 == io_inputs_1 ? 7'h0 : _GEN_3672; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3674 = 10'h15a == io_inputs_1 ? 7'h0 : _GEN_3673; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3675 = 10'h15b == io_inputs_1 ? 7'h0 : _GEN_3674; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3676 = 10'h15c == io_inputs_1 ? 7'h0 : _GEN_3675; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3677 = 10'h15d == io_inputs_1 ? 7'h0 : _GEN_3676; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3678 = 10'h15e == io_inputs_1 ? 7'h0 : _GEN_3677; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3679 = 10'h15f == io_inputs_1 ? 7'h0 : _GEN_3678; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3680 = 10'h160 == io_inputs_1 ? 7'h0 : _GEN_3679; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3681 = 10'h161 == io_inputs_1 ? 7'h0 : _GEN_3680; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3682 = 10'h162 == io_inputs_1 ? 7'h0 : _GEN_3681; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3683 = 10'h163 == io_inputs_1 ? 7'h0 : _GEN_3682; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3684 = 10'h164 == io_inputs_1 ? 7'h0 : _GEN_3683; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3685 = 10'h165 == io_inputs_1 ? 7'h0 : _GEN_3684; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3686 = 10'h166 == io_inputs_1 ? 7'h0 : _GEN_3685; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3687 = 10'h167 == io_inputs_1 ? 7'h0 : _GEN_3686; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3688 = 10'h168 == io_inputs_1 ? 7'h0 : _GEN_3687; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3689 = 10'h169 == io_inputs_1 ? 7'h0 : _GEN_3688; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3690 = 10'h16a == io_inputs_1 ? 7'h0 : _GEN_3689; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3691 = 10'h16b == io_inputs_1 ? 7'h0 : _GEN_3690; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3692 = 10'h16c == io_inputs_1 ? 7'h0 : _GEN_3691; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3693 = 10'h16d == io_inputs_1 ? 7'h0 : _GEN_3692; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3694 = 10'h16e == io_inputs_1 ? 7'h0 : _GEN_3693; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3695 = 10'h16f == io_inputs_1 ? 7'h0 : _GEN_3694; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3696 = 10'h170 == io_inputs_1 ? 7'h0 : _GEN_3695; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3697 = 10'h171 == io_inputs_1 ? 7'h0 : _GEN_3696; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3698 = 10'h172 == io_inputs_1 ? 7'h0 : _GEN_3697; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3699 = 10'h173 == io_inputs_1 ? 7'h0 : _GEN_3698; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3700 = 10'h174 == io_inputs_1 ? 7'h0 : _GEN_3699; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3701 = 10'h175 == io_inputs_1 ? 7'h0 : _GEN_3700; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3702 = 10'h176 == io_inputs_1 ? 7'h0 : _GEN_3701; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3703 = 10'h177 == io_inputs_1 ? 7'h0 : _GEN_3702; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3704 = 10'h178 == io_inputs_1 ? 7'h0 : _GEN_3703; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3705 = 10'h179 == io_inputs_1 ? 7'h0 : _GEN_3704; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3706 = 10'h17a == io_inputs_1 ? 7'h0 : _GEN_3705; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3707 = 10'h17b == io_inputs_1 ? 7'h0 : _GEN_3706; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3708 = 10'h17c == io_inputs_1 ? 7'h0 : _GEN_3707; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3709 = 10'h17d == io_inputs_1 ? 7'h0 : _GEN_3708; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3710 = 10'h17e == io_inputs_1 ? 7'h0 : _GEN_3709; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3711 = 10'h17f == io_inputs_1 ? 7'h0 : _GEN_3710; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3712 = 10'h180 == io_inputs_1 ? 7'h0 : _GEN_3711; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3713 = 10'h181 == io_inputs_1 ? 7'h0 : _GEN_3712; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3714 = 10'h182 == io_inputs_1 ? 7'h0 : _GEN_3713; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3715 = 10'h183 == io_inputs_1 ? 7'h0 : _GEN_3714; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3716 = 10'h184 == io_inputs_1 ? 7'h0 : _GEN_3715; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3717 = 10'h185 == io_inputs_1 ? 7'h0 : _GEN_3716; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3718 = 10'h186 == io_inputs_1 ? 7'h0 : _GEN_3717; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3719 = 10'h187 == io_inputs_1 ? 7'h0 : _GEN_3718; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3720 = 10'h188 == io_inputs_1 ? 7'h0 : _GEN_3719; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3721 = 10'h189 == io_inputs_1 ? 7'h0 : _GEN_3720; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3722 = 10'h18a == io_inputs_1 ? 7'h0 : _GEN_3721; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3723 = 10'h18b == io_inputs_1 ? 7'h0 : _GEN_3722; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3724 = 10'h18c == io_inputs_1 ? 7'h0 : _GEN_3723; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3725 = 10'h18d == io_inputs_1 ? 7'h0 : _GEN_3724; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3726 = 10'h18e == io_inputs_1 ? 7'h0 : _GEN_3725; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3727 = 10'h18f == io_inputs_1 ? 7'h0 : _GEN_3726; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3728 = 10'h190 == io_inputs_1 ? 7'h0 : _GEN_3727; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3729 = 10'h191 == io_inputs_1 ? 7'h0 : _GEN_3728; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3730 = 10'h192 == io_inputs_1 ? 7'h0 : _GEN_3729; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3731 = 10'h193 == io_inputs_1 ? 7'h0 : _GEN_3730; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3732 = 10'h194 == io_inputs_1 ? 7'h0 : _GEN_3731; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3733 = 10'h195 == io_inputs_1 ? 7'h0 : _GEN_3732; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3734 = 10'h196 == io_inputs_1 ? 7'h0 : _GEN_3733; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3735 = 10'h197 == io_inputs_1 ? 7'h0 : _GEN_3734; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3736 = 10'h198 == io_inputs_1 ? 7'h0 : _GEN_3735; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3737 = 10'h199 == io_inputs_1 ? 7'h0 : _GEN_3736; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3738 = 10'h19a == io_inputs_1 ? 7'h0 : _GEN_3737; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3739 = 10'h19b == io_inputs_1 ? 7'h0 : _GEN_3738; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3740 = 10'h19c == io_inputs_1 ? 7'h0 : _GEN_3739; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3741 = 10'h19d == io_inputs_1 ? 7'h0 : _GEN_3740; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3742 = 10'h19e == io_inputs_1 ? 7'h0 : _GEN_3741; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3743 = 10'h19f == io_inputs_1 ? 7'h0 : _GEN_3742; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3744 = 10'h1a0 == io_inputs_1 ? 7'h0 : _GEN_3743; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3745 = 10'h1a1 == io_inputs_1 ? 7'h0 : _GEN_3744; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3746 = 10'h1a2 == io_inputs_1 ? 7'h0 : _GEN_3745; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3747 = 10'h1a3 == io_inputs_1 ? 7'h0 : _GEN_3746; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3748 = 10'h1a4 == io_inputs_1 ? 7'h0 : _GEN_3747; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3749 = 10'h1a5 == io_inputs_1 ? 7'h0 : _GEN_3748; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3750 = 10'h1a6 == io_inputs_1 ? 7'h0 : _GEN_3749; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3751 = 10'h1a7 == io_inputs_1 ? 7'h0 : _GEN_3750; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3752 = 10'h1a8 == io_inputs_1 ? 7'h0 : _GEN_3751; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3753 = 10'h1a9 == io_inputs_1 ? 7'h0 : _GEN_3752; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3754 = 10'h1aa == io_inputs_1 ? 7'h0 : _GEN_3753; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3755 = 10'h1ab == io_inputs_1 ? 7'h0 : _GEN_3754; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3756 = 10'h1ac == io_inputs_1 ? 7'h0 : _GEN_3755; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3757 = 10'h1ad == io_inputs_1 ? 7'h0 : _GEN_3756; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3758 = 10'h1ae == io_inputs_1 ? 7'h0 : _GEN_3757; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3759 = 10'h1af == io_inputs_1 ? 7'h0 : _GEN_3758; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3760 = 10'h1b0 == io_inputs_1 ? 7'h0 : _GEN_3759; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3761 = 10'h1b1 == io_inputs_1 ? 7'h0 : _GEN_3760; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3762 = 10'h1b2 == io_inputs_1 ? 7'h0 : _GEN_3761; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3763 = 10'h1b3 == io_inputs_1 ? 7'h0 : _GEN_3762; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3764 = 10'h1b4 == io_inputs_1 ? 7'h0 : _GEN_3763; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3765 = 10'h1b5 == io_inputs_1 ? 7'h0 : _GEN_3764; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3766 = 10'h1b6 == io_inputs_1 ? 7'h0 : _GEN_3765; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3767 = 10'h1b7 == io_inputs_1 ? 7'h0 : _GEN_3766; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3768 = 10'h1b8 == io_inputs_1 ? 7'h0 : _GEN_3767; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3769 = 10'h1b9 == io_inputs_1 ? 7'h0 : _GEN_3768; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3770 = 10'h1ba == io_inputs_1 ? 7'h0 : _GEN_3769; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3771 = 10'h1bb == io_inputs_1 ? 7'h0 : _GEN_3770; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3772 = 10'h1bc == io_inputs_1 ? 7'h0 : _GEN_3771; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3773 = 10'h1bd == io_inputs_1 ? 7'h0 : _GEN_3772; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3774 = 10'h1be == io_inputs_1 ? 7'h0 : _GEN_3773; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3775 = 10'h1bf == io_inputs_1 ? 7'h0 : _GEN_3774; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3776 = 10'h1c0 == io_inputs_1 ? 7'h0 : _GEN_3775; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3777 = 10'h1c1 == io_inputs_1 ? 7'h0 : _GEN_3776; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3778 = 10'h1c2 == io_inputs_1 ? 7'h0 : _GEN_3777; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3779 = 10'h1c3 == io_inputs_1 ? 7'h0 : _GEN_3778; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3780 = 10'h1c4 == io_inputs_1 ? 7'h0 : _GEN_3779; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3781 = 10'h1c5 == io_inputs_1 ? 7'h0 : _GEN_3780; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3782 = 10'h1c6 == io_inputs_1 ? 7'h0 : _GEN_3781; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3783 = 10'h1c7 == io_inputs_1 ? 7'h0 : _GEN_3782; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3784 = 10'h1c8 == io_inputs_1 ? 7'h0 : _GEN_3783; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3785 = 10'h1c9 == io_inputs_1 ? 7'h0 : _GEN_3784; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3786 = 10'h1ca == io_inputs_1 ? 7'h0 : _GEN_3785; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3787 = 10'h1cb == io_inputs_1 ? 7'h0 : _GEN_3786; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3788 = 10'h1cc == io_inputs_1 ? 7'h0 : _GEN_3787; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3789 = 10'h1cd == io_inputs_1 ? 7'h0 : _GEN_3788; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3790 = 10'h1ce == io_inputs_1 ? 7'h0 : _GEN_3789; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3791 = 10'h1cf == io_inputs_1 ? 7'h0 : _GEN_3790; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3792 = 10'h1d0 == io_inputs_1 ? 7'h0 : _GEN_3791; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3793 = 10'h1d1 == io_inputs_1 ? 7'h0 : _GEN_3792; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3794 = 10'h1d2 == io_inputs_1 ? 7'h0 : _GEN_3793; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3795 = 10'h1d3 == io_inputs_1 ? 7'h0 : _GEN_3794; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3796 = 10'h1d4 == io_inputs_1 ? 7'h0 : _GEN_3795; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3797 = 10'h1d5 == io_inputs_1 ? 7'h0 : _GEN_3796; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3798 = 10'h1d6 == io_inputs_1 ? 7'h0 : _GEN_3797; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3799 = 10'h1d7 == io_inputs_1 ? 7'h0 : _GEN_3798; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3800 = 10'h1d8 == io_inputs_1 ? 7'h0 : _GEN_3799; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3801 = 10'h1d9 == io_inputs_1 ? 7'h0 : _GEN_3800; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3802 = 10'h1da == io_inputs_1 ? 7'h0 : _GEN_3801; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3803 = 10'h1db == io_inputs_1 ? 7'h0 : _GEN_3802; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3804 = 10'h1dc == io_inputs_1 ? 7'h0 : _GEN_3803; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3805 = 10'h1dd == io_inputs_1 ? 7'h0 : _GEN_3804; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3806 = 10'h1de == io_inputs_1 ? 7'h0 : _GEN_3805; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3807 = 10'h1df == io_inputs_1 ? 7'h0 : _GEN_3806; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3808 = 10'h1e0 == io_inputs_1 ? 7'h0 : _GEN_3807; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3809 = 10'h1e1 == io_inputs_1 ? 7'h0 : _GEN_3808; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3810 = 10'h1e2 == io_inputs_1 ? 7'h0 : _GEN_3809; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3811 = 10'h1e3 == io_inputs_1 ? 7'h0 : _GEN_3810; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3812 = 10'h1e4 == io_inputs_1 ? 7'h0 : _GEN_3811; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3813 = 10'h1e5 == io_inputs_1 ? 7'h0 : _GEN_3812; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3814 = 10'h1e6 == io_inputs_1 ? 7'h0 : _GEN_3813; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3815 = 10'h1e7 == io_inputs_1 ? 7'h0 : _GEN_3814; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3816 = 10'h1e8 == io_inputs_1 ? 7'h0 : _GEN_3815; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3817 = 10'h1e9 == io_inputs_1 ? 7'h0 : _GEN_3816; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3818 = 10'h1ea == io_inputs_1 ? 7'h0 : _GEN_3817; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3819 = 10'h1eb == io_inputs_1 ? 7'h0 : _GEN_3818; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3820 = 10'h1ec == io_inputs_1 ? 7'h0 : _GEN_3819; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3821 = 10'h1ed == io_inputs_1 ? 7'h0 : _GEN_3820; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3822 = 10'h1ee == io_inputs_1 ? 7'h0 : _GEN_3821; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3823 = 10'h1ef == io_inputs_1 ? 7'h0 : _GEN_3822; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3824 = 10'h1f0 == io_inputs_1 ? 7'h0 : _GEN_3823; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3825 = 10'h1f1 == io_inputs_1 ? 7'h0 : _GEN_3824; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3826 = 10'h1f2 == io_inputs_1 ? 7'h0 : _GEN_3825; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3827 = 10'h1f3 == io_inputs_1 ? 7'h0 : _GEN_3826; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3828 = 10'h1f4 == io_inputs_1 ? 7'h0 : _GEN_3827; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3829 = 10'h1f5 == io_inputs_1 ? 7'h0 : _GEN_3828; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3830 = 10'h1f6 == io_inputs_1 ? 7'h0 : _GEN_3829; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3831 = 10'h1f7 == io_inputs_1 ? 7'h0 : _GEN_3830; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3832 = 10'h1f8 == io_inputs_1 ? 7'h0 : _GEN_3831; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3833 = 10'h1f9 == io_inputs_1 ? 7'h0 : _GEN_3832; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3834 = 10'h1fa == io_inputs_1 ? 7'h0 : _GEN_3833; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3835 = 10'h1fb == io_inputs_1 ? 7'h0 : _GEN_3834; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3836 = 10'h1fc == io_inputs_1 ? 7'h0 : _GEN_3835; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3837 = 10'h1fd == io_inputs_1 ? 7'h0 : _GEN_3836; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3838 = 10'h1fe == io_inputs_1 ? 7'h0 : _GEN_3837; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3839 = 10'h1ff == io_inputs_1 ? 7'h0 : _GEN_3838; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3840 = 10'h200 == io_inputs_1 ? 7'h0 : _GEN_3839; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3841 = 10'h201 == io_inputs_1 ? 7'h0 : _GEN_3840; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3842 = 10'h202 == io_inputs_1 ? 7'h0 : _GEN_3841; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3843 = 10'h203 == io_inputs_1 ? 7'h0 : _GEN_3842; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3844 = 10'h204 == io_inputs_1 ? 7'h0 : _GEN_3843; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3845 = 10'h205 == io_inputs_1 ? 7'h0 : _GEN_3844; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3846 = 10'h206 == io_inputs_1 ? 7'h0 : _GEN_3845; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3847 = 10'h207 == io_inputs_1 ? 7'h0 : _GEN_3846; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3848 = 10'h208 == io_inputs_1 ? 7'h0 : _GEN_3847; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3849 = 10'h209 == io_inputs_1 ? 7'h0 : _GEN_3848; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3850 = 10'h20a == io_inputs_1 ? 7'h0 : _GEN_3849; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3851 = 10'h20b == io_inputs_1 ? 7'h0 : _GEN_3850; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3852 = 10'h20c == io_inputs_1 ? 7'h0 : _GEN_3851; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3853 = 10'h20d == io_inputs_1 ? 7'h0 : _GEN_3852; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3854 = 10'h20e == io_inputs_1 ? 7'h0 : _GEN_3853; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3855 = 10'h20f == io_inputs_1 ? 7'h0 : _GEN_3854; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3856 = 10'h210 == io_inputs_1 ? 7'h0 : _GEN_3855; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3857 = 10'h211 == io_inputs_1 ? 7'h0 : _GEN_3856; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3858 = 10'h212 == io_inputs_1 ? 7'h0 : _GEN_3857; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3859 = 10'h213 == io_inputs_1 ? 7'h0 : _GEN_3858; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3860 = 10'h214 == io_inputs_1 ? 7'h0 : _GEN_3859; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3861 = 10'h215 == io_inputs_1 ? 7'h0 : _GEN_3860; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3862 = 10'h216 == io_inputs_1 ? 7'h0 : _GEN_3861; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3863 = 10'h217 == io_inputs_1 ? 7'h0 : _GEN_3862; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3864 = 10'h218 == io_inputs_1 ? 7'h0 : _GEN_3863; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3865 = 10'h219 == io_inputs_1 ? 7'h0 : _GEN_3864; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3866 = 10'h21a == io_inputs_1 ? 7'h0 : _GEN_3865; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3867 = 10'h21b == io_inputs_1 ? 7'h0 : _GEN_3866; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3868 = 10'h21c == io_inputs_1 ? 7'h0 : _GEN_3867; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3869 = 10'h21d == io_inputs_1 ? 7'h0 : _GEN_3868; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3870 = 10'h21e == io_inputs_1 ? 7'h0 : _GEN_3869; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3871 = 10'h21f == io_inputs_1 ? 7'h0 : _GEN_3870; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3872 = 10'h220 == io_inputs_1 ? 7'h0 : _GEN_3871; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3873 = 10'h221 == io_inputs_1 ? 7'h0 : _GEN_3872; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3874 = 10'h222 == io_inputs_1 ? 7'h0 : _GEN_3873; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3875 = 10'h223 == io_inputs_1 ? 7'h0 : _GEN_3874; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3876 = 10'h224 == io_inputs_1 ? 7'h0 : _GEN_3875; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3877 = 10'h225 == io_inputs_1 ? 7'h0 : _GEN_3876; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3878 = 10'h226 == io_inputs_1 ? 7'h0 : _GEN_3877; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3879 = 10'h227 == io_inputs_1 ? 7'h0 : _GEN_3878; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3880 = 10'h228 == io_inputs_1 ? 7'h0 : _GEN_3879; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3881 = 10'h229 == io_inputs_1 ? 7'h0 : _GEN_3880; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3882 = 10'h22a == io_inputs_1 ? 7'h0 : _GEN_3881; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3883 = 10'h22b == io_inputs_1 ? 7'h0 : _GEN_3882; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3884 = 10'h22c == io_inputs_1 ? 7'h0 : _GEN_3883; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3885 = 10'h22d == io_inputs_1 ? 7'h0 : _GEN_3884; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3886 = 10'h22e == io_inputs_1 ? 7'h0 : _GEN_3885; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3887 = 10'h22f == io_inputs_1 ? 7'h0 : _GEN_3886; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3888 = 10'h230 == io_inputs_1 ? 7'h0 : _GEN_3887; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3889 = 10'h231 == io_inputs_1 ? 7'h0 : _GEN_3888; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3890 = 10'h232 == io_inputs_1 ? 7'h0 : _GEN_3889; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3891 = 10'h233 == io_inputs_1 ? 7'h0 : _GEN_3890; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3892 = 10'h234 == io_inputs_1 ? 7'h0 : _GEN_3891; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3893 = 10'h235 == io_inputs_1 ? 7'h0 : _GEN_3892; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3894 = 10'h236 == io_inputs_1 ? 7'h0 : _GEN_3893; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3895 = 10'h237 == io_inputs_1 ? 7'h0 : _GEN_3894; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3896 = 10'h238 == io_inputs_1 ? 7'h0 : _GEN_3895; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3897 = 10'h239 == io_inputs_1 ? 7'h0 : _GEN_3896; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3898 = 10'h23a == io_inputs_1 ? 7'h0 : _GEN_3897; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3899 = 10'h23b == io_inputs_1 ? 7'h0 : _GEN_3898; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3900 = 10'h23c == io_inputs_1 ? 7'h0 : _GEN_3899; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3901 = 10'h23d == io_inputs_1 ? 7'h0 : _GEN_3900; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3902 = 10'h23e == io_inputs_1 ? 7'h0 : _GEN_3901; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3903 = 10'h23f == io_inputs_1 ? 7'h0 : _GEN_3902; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3904 = 10'h240 == io_inputs_1 ? 7'h0 : _GEN_3903; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3905 = 10'h241 == io_inputs_1 ? 7'h0 : _GEN_3904; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3906 = 10'h242 == io_inputs_1 ? 7'h0 : _GEN_3905; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3907 = 10'h243 == io_inputs_1 ? 7'h0 : _GEN_3906; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3908 = 10'h244 == io_inputs_1 ? 7'h0 : _GEN_3907; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3909 = 10'h245 == io_inputs_1 ? 7'h0 : _GEN_3908; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3910 = 10'h246 == io_inputs_1 ? 7'h0 : _GEN_3909; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3911 = 10'h247 == io_inputs_1 ? 7'h0 : _GEN_3910; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3912 = 10'h248 == io_inputs_1 ? 7'h0 : _GEN_3911; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3913 = 10'h249 == io_inputs_1 ? 7'h0 : _GEN_3912; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3914 = 10'h24a == io_inputs_1 ? 7'h0 : _GEN_3913; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3915 = 10'h24b == io_inputs_1 ? 7'h0 : _GEN_3914; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3916 = 10'h24c == io_inputs_1 ? 7'h0 : _GEN_3915; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3917 = 10'h24d == io_inputs_1 ? 7'h0 : _GEN_3916; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3918 = 10'h24e == io_inputs_1 ? 7'h0 : _GEN_3917; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3919 = 10'h24f == io_inputs_1 ? 7'h0 : _GEN_3918; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3920 = 10'h250 == io_inputs_1 ? 7'h0 : _GEN_3919; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3921 = 10'h251 == io_inputs_1 ? 7'h0 : _GEN_3920; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3922 = 10'h252 == io_inputs_1 ? 7'h0 : _GEN_3921; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3923 = 10'h253 == io_inputs_1 ? 7'h0 : _GEN_3922; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3924 = 10'h254 == io_inputs_1 ? 7'h0 : _GEN_3923; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3925 = 10'h255 == io_inputs_1 ? 7'h0 : _GEN_3924; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3926 = 10'h256 == io_inputs_1 ? 7'h0 : _GEN_3925; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3927 = 10'h257 == io_inputs_1 ? 7'h0 : _GEN_3926; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3928 = 10'h258 == io_inputs_1 ? 7'h0 : _GEN_3927; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3929 = 10'h259 == io_inputs_1 ? 7'h0 : _GEN_3928; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3930 = 10'h25a == io_inputs_1 ? 7'h0 : _GEN_3929; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3931 = 10'h25b == io_inputs_1 ? 7'h0 : _GEN_3930; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3932 = 10'h25c == io_inputs_1 ? 7'h0 : _GEN_3931; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3933 = 10'h25d == io_inputs_1 ? 7'h0 : _GEN_3932; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3934 = 10'h25e == io_inputs_1 ? 7'h0 : _GEN_3933; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3935 = 10'h25f == io_inputs_1 ? 7'h0 : _GEN_3934; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3936 = 10'h260 == io_inputs_1 ? 7'h0 : _GEN_3935; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3937 = 10'h261 == io_inputs_1 ? 7'h0 : _GEN_3936; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3938 = 10'h262 == io_inputs_1 ? 7'h0 : _GEN_3937; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3939 = 10'h263 == io_inputs_1 ? 7'h0 : _GEN_3938; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3940 = 10'h264 == io_inputs_1 ? 7'h0 : _GEN_3939; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3941 = 10'h265 == io_inputs_1 ? 7'h0 : _GEN_3940; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3942 = 10'h266 == io_inputs_1 ? 7'h0 : _GEN_3941; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3943 = 10'h267 == io_inputs_1 ? 7'h0 : _GEN_3942; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3944 = 10'h268 == io_inputs_1 ? 7'h0 : _GEN_3943; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3945 = 10'h269 == io_inputs_1 ? 7'h0 : _GEN_3944; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3946 = 10'h26a == io_inputs_1 ? 7'h0 : _GEN_3945; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3947 = 10'h26b == io_inputs_1 ? 7'h0 : _GEN_3946; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3948 = 10'h26c == io_inputs_1 ? 7'h0 : _GEN_3947; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3949 = 10'h26d == io_inputs_1 ? 7'h0 : _GEN_3948; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3950 = 10'h26e == io_inputs_1 ? 7'h0 : _GEN_3949; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3951 = 10'h26f == io_inputs_1 ? 7'h0 : _GEN_3950; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3952 = 10'h270 == io_inputs_1 ? 7'h0 : _GEN_3951; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3953 = 10'h271 == io_inputs_1 ? 7'h0 : _GEN_3952; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3954 = 10'h272 == io_inputs_1 ? 7'h0 : _GEN_3953; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3955 = 10'h273 == io_inputs_1 ? 7'h0 : _GEN_3954; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3956 = 10'h274 == io_inputs_1 ? 7'h0 : _GEN_3955; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3957 = 10'h275 == io_inputs_1 ? 7'h0 : _GEN_3956; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3958 = 10'h276 == io_inputs_1 ? 7'h0 : _GEN_3957; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3959 = 10'h277 == io_inputs_1 ? 7'h0 : _GEN_3958; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3960 = 10'h278 == io_inputs_1 ? 7'h0 : _GEN_3959; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3961 = 10'h279 == io_inputs_1 ? 7'h0 : _GEN_3960; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3962 = 10'h27a == io_inputs_1 ? 7'h0 : _GEN_3961; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3963 = 10'h27b == io_inputs_1 ? 7'h0 : _GEN_3962; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3964 = 10'h27c == io_inputs_1 ? 7'h0 : _GEN_3963; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3965 = 10'h27d == io_inputs_1 ? 7'h0 : _GEN_3964; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3966 = 10'h27e == io_inputs_1 ? 7'h0 : _GEN_3965; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3967 = 10'h27f == io_inputs_1 ? 7'h0 : _GEN_3966; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3968 = 10'h280 == io_inputs_1 ? 7'h0 : _GEN_3967; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3969 = 10'h281 == io_inputs_1 ? 7'h0 : _GEN_3968; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3970 = 10'h282 == io_inputs_1 ? 7'h0 : _GEN_3969; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3971 = 10'h283 == io_inputs_1 ? 7'h0 : _GEN_3970; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3972 = 10'h284 == io_inputs_1 ? 7'h0 : _GEN_3971; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3973 = 10'h285 == io_inputs_1 ? 7'h0 : _GEN_3972; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3974 = 10'h286 == io_inputs_1 ? 7'h0 : _GEN_3973; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3975 = 10'h287 == io_inputs_1 ? 7'h0 : _GEN_3974; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3976 = 10'h288 == io_inputs_1 ? 7'h0 : _GEN_3975; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3977 = 10'h289 == io_inputs_1 ? 7'h0 : _GEN_3976; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3978 = 10'h28a == io_inputs_1 ? 7'h0 : _GEN_3977; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3979 = 10'h28b == io_inputs_1 ? 7'h0 : _GEN_3978; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3980 = 10'h28c == io_inputs_1 ? 7'h0 : _GEN_3979; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3981 = 10'h28d == io_inputs_1 ? 7'h0 : _GEN_3980; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3982 = 10'h28e == io_inputs_1 ? 7'h0 : _GEN_3981; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3983 = 10'h28f == io_inputs_1 ? 7'h0 : _GEN_3982; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3984 = 10'h290 == io_inputs_1 ? 7'h0 : _GEN_3983; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3985 = 10'h291 == io_inputs_1 ? 7'h0 : _GEN_3984; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3986 = 10'h292 == io_inputs_1 ? 7'h0 : _GEN_3985; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3987 = 10'h293 == io_inputs_1 ? 7'h0 : _GEN_3986; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3988 = 10'h294 == io_inputs_1 ? 7'h0 : _GEN_3987; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3989 = 10'h295 == io_inputs_1 ? 7'h0 : _GEN_3988; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3990 = 10'h296 == io_inputs_1 ? 7'h0 : _GEN_3989; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3991 = 10'h297 == io_inputs_1 ? 7'h0 : _GEN_3990; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3992 = 10'h298 == io_inputs_1 ? 7'h0 : _GEN_3991; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3993 = 10'h299 == io_inputs_1 ? 7'h0 : _GEN_3992; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3994 = 10'h29a == io_inputs_1 ? 7'h0 : _GEN_3993; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3995 = 10'h29b == io_inputs_1 ? 7'h0 : _GEN_3994; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3996 = 10'h29c == io_inputs_1 ? 7'h0 : _GEN_3995; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3997 = 10'h29d == io_inputs_1 ? 7'h0 : _GEN_3996; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3998 = 10'h29e == io_inputs_1 ? 7'h0 : _GEN_3997; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_3999 = 10'h29f == io_inputs_1 ? 7'h0 : _GEN_3998; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4000 = 10'h2a0 == io_inputs_1 ? 7'h0 : _GEN_3999; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4001 = 10'h2a1 == io_inputs_1 ? 7'h0 : _GEN_4000; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4002 = 10'h2a2 == io_inputs_1 ? 7'h0 : _GEN_4001; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4003 = 10'h2a3 == io_inputs_1 ? 7'h0 : _GEN_4002; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4004 = 10'h2a4 == io_inputs_1 ? 7'h0 : _GEN_4003; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4005 = 10'h2a5 == io_inputs_1 ? 7'h0 : _GEN_4004; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4006 = 10'h2a6 == io_inputs_1 ? 7'h0 : _GEN_4005; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4007 = 10'h2a7 == io_inputs_1 ? 7'h0 : _GEN_4006; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4008 = 10'h2a8 == io_inputs_1 ? 7'h0 : _GEN_4007; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4009 = 10'h2a9 == io_inputs_1 ? 7'h0 : _GEN_4008; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4010 = 10'h2aa == io_inputs_1 ? 7'h0 : _GEN_4009; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4011 = 10'h2ab == io_inputs_1 ? 7'h0 : _GEN_4010; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4012 = 10'h2ac == io_inputs_1 ? 7'h0 : _GEN_4011; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4013 = 10'h2ad == io_inputs_1 ? 7'h0 : _GEN_4012; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4014 = 10'h2ae == io_inputs_1 ? 7'h0 : _GEN_4013; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4015 = 10'h2af == io_inputs_1 ? 7'h0 : _GEN_4014; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4016 = 10'h2b0 == io_inputs_1 ? 7'h0 : _GEN_4015; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4017 = 10'h2b1 == io_inputs_1 ? 7'h0 : _GEN_4016; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4018 = 10'h2b2 == io_inputs_1 ? 7'h0 : _GEN_4017; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4019 = 10'h2b3 == io_inputs_1 ? 7'h0 : _GEN_4018; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4020 = 10'h2b4 == io_inputs_1 ? 7'h0 : _GEN_4019; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4021 = 10'h2b5 == io_inputs_1 ? 7'h0 : _GEN_4020; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4022 = 10'h2b6 == io_inputs_1 ? 7'h0 : _GEN_4021; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4023 = 10'h2b7 == io_inputs_1 ? 7'h0 : _GEN_4022; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4024 = 10'h2b8 == io_inputs_1 ? 7'h0 : _GEN_4023; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4025 = 10'h2b9 == io_inputs_1 ? 7'h0 : _GEN_4024; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4026 = 10'h2ba == io_inputs_1 ? 7'h0 : _GEN_4025; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4027 = 10'h2bb == io_inputs_1 ? 7'h0 : _GEN_4026; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4028 = 10'h2bc == io_inputs_1 ? 7'h0 : _GEN_4027; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4029 = 10'h2bd == io_inputs_1 ? 7'h0 : _GEN_4028; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4030 = 10'h2be == io_inputs_1 ? 7'h0 : _GEN_4029; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4031 = 10'h2bf == io_inputs_1 ? 7'h0 : _GEN_4030; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4032 = 10'h2c0 == io_inputs_1 ? 7'h0 : _GEN_4031; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4033 = 10'h2c1 == io_inputs_1 ? 7'h0 : _GEN_4032; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4034 = 10'h2c2 == io_inputs_1 ? 7'h0 : _GEN_4033; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4035 = 10'h2c3 == io_inputs_1 ? 7'h0 : _GEN_4034; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4036 = 10'h2c4 == io_inputs_1 ? 7'h0 : _GEN_4035; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4037 = 10'h2c5 == io_inputs_1 ? 7'h0 : _GEN_4036; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4038 = 10'h2c6 == io_inputs_1 ? 7'h0 : _GEN_4037; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4039 = 10'h2c7 == io_inputs_1 ? 7'h0 : _GEN_4038; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4040 = 10'h2c8 == io_inputs_1 ? 7'h0 : _GEN_4039; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4041 = 10'h2c9 == io_inputs_1 ? 7'h0 : _GEN_4040; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4042 = 10'h2ca == io_inputs_1 ? 7'h0 : _GEN_4041; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4043 = 10'h2cb == io_inputs_1 ? 7'h0 : _GEN_4042; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4044 = 10'h2cc == io_inputs_1 ? 7'h0 : _GEN_4043; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4045 = 10'h2cd == io_inputs_1 ? 7'h0 : _GEN_4044; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4046 = 10'h2ce == io_inputs_1 ? 7'h0 : _GEN_4045; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4047 = 10'h2cf == io_inputs_1 ? 7'h0 : _GEN_4046; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4048 = 10'h2d0 == io_inputs_1 ? 7'h0 : _GEN_4047; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4049 = 10'h2d1 == io_inputs_1 ? 7'h0 : _GEN_4048; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4050 = 10'h2d2 == io_inputs_1 ? 7'h0 : _GEN_4049; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4051 = 10'h2d3 == io_inputs_1 ? 7'h0 : _GEN_4050; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4052 = 10'h2d4 == io_inputs_1 ? 7'h0 : _GEN_4051; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4053 = 10'h2d5 == io_inputs_1 ? 7'h0 : _GEN_4052; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4054 = 10'h2d6 == io_inputs_1 ? 7'h0 : _GEN_4053; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4055 = 10'h2d7 == io_inputs_1 ? 7'h0 : _GEN_4054; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4056 = 10'h2d8 == io_inputs_1 ? 7'h0 : _GEN_4055; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4057 = 10'h2d9 == io_inputs_1 ? 7'h0 : _GEN_4056; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4058 = 10'h2da == io_inputs_1 ? 7'h0 : _GEN_4057; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4059 = 10'h2db == io_inputs_1 ? 7'h0 : _GEN_4058; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4060 = 10'h2dc == io_inputs_1 ? 7'h0 : _GEN_4059; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4061 = 10'h2dd == io_inputs_1 ? 7'h0 : _GEN_4060; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4062 = 10'h2de == io_inputs_1 ? 7'h0 : _GEN_4061; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4063 = 10'h2df == io_inputs_1 ? 7'h0 : _GEN_4062; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4064 = 10'h2e0 == io_inputs_1 ? 7'h0 : _GEN_4063; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4065 = 10'h2e1 == io_inputs_1 ? 7'h0 : _GEN_4064; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4066 = 10'h2e2 == io_inputs_1 ? 7'h0 : _GEN_4065; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4067 = 10'h2e3 == io_inputs_1 ? 7'h0 : _GEN_4066; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4068 = 10'h2e4 == io_inputs_1 ? 7'h0 : _GEN_4067; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4069 = 10'h2e5 == io_inputs_1 ? 7'h0 : _GEN_4068; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4070 = 10'h2e6 == io_inputs_1 ? 7'h0 : _GEN_4069; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4071 = 10'h2e7 == io_inputs_1 ? 7'h0 : _GEN_4070; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4072 = 10'h2e8 == io_inputs_1 ? 7'h0 : _GEN_4071; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4073 = 10'h2e9 == io_inputs_1 ? 7'h0 : _GEN_4072; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4074 = 10'h2ea == io_inputs_1 ? 7'h0 : _GEN_4073; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4075 = 10'h2eb == io_inputs_1 ? 7'h0 : _GEN_4074; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4076 = 10'h2ec == io_inputs_1 ? 7'h0 : _GEN_4075; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4077 = 10'h2ed == io_inputs_1 ? 7'h0 : _GEN_4076; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4078 = 10'h2ee == io_inputs_1 ? 7'h0 : _GEN_4077; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4079 = 10'h2ef == io_inputs_1 ? 7'h0 : _GEN_4078; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4080 = 10'h2f0 == io_inputs_1 ? 7'h0 : _GEN_4079; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4081 = 10'h2f1 == io_inputs_1 ? 7'h0 : _GEN_4080; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4082 = 10'h2f2 == io_inputs_1 ? 7'h0 : _GEN_4081; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4083 = 10'h2f3 == io_inputs_1 ? 7'h0 : _GEN_4082; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4084 = 10'h2f4 == io_inputs_1 ? 7'h0 : _GEN_4083; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4085 = 10'h2f5 == io_inputs_1 ? 7'h0 : _GEN_4084; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4086 = 10'h2f6 == io_inputs_1 ? 7'h0 : _GEN_4085; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4087 = 10'h2f7 == io_inputs_1 ? 7'h0 : _GEN_4086; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4088 = 10'h2f8 == io_inputs_1 ? 7'h0 : _GEN_4087; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4089 = 10'h2f9 == io_inputs_1 ? 7'h0 : _GEN_4088; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4090 = 10'h2fa == io_inputs_1 ? 7'h0 : _GEN_4089; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4091 = 10'h2fb == io_inputs_1 ? 7'h0 : _GEN_4090; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4092 = 10'h2fc == io_inputs_1 ? 7'h0 : _GEN_4091; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4093 = 10'h2fd == io_inputs_1 ? 7'h0 : _GEN_4092; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4094 = 10'h2fe == io_inputs_1 ? 7'h0 : _GEN_4093; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4095 = 10'h2ff == io_inputs_1 ? 7'h0 : _GEN_4094; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4096 = 10'h300 == io_inputs_1 ? 7'h0 : _GEN_4095; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4097 = 10'h301 == io_inputs_1 ? 7'h0 : _GEN_4096; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4098 = 10'h302 == io_inputs_1 ? 7'h0 : _GEN_4097; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4099 = 10'h303 == io_inputs_1 ? 7'h0 : _GEN_4098; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4100 = 10'h304 == io_inputs_1 ? 7'h0 : _GEN_4099; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4101 = 10'h305 == io_inputs_1 ? 7'h0 : _GEN_4100; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4102 = 10'h306 == io_inputs_1 ? 7'h0 : _GEN_4101; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4103 = 10'h307 == io_inputs_1 ? 7'h0 : _GEN_4102; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4104 = 10'h308 == io_inputs_1 ? 7'h0 : _GEN_4103; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4105 = 10'h309 == io_inputs_1 ? 7'h0 : _GEN_4104; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4106 = 10'h30a == io_inputs_1 ? 7'h0 : _GEN_4105; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4107 = 10'h30b == io_inputs_1 ? 7'h0 : _GEN_4106; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4108 = 10'h30c == io_inputs_1 ? 7'h0 : _GEN_4107; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4109 = 10'h30d == io_inputs_1 ? 7'h0 : _GEN_4108; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4110 = 10'h30e == io_inputs_1 ? 7'h0 : _GEN_4109; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4111 = 10'h30f == io_inputs_1 ? 7'h0 : _GEN_4110; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4112 = 10'h310 == io_inputs_1 ? 7'h0 : _GEN_4111; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4113 = 10'h311 == io_inputs_1 ? 7'h0 : _GEN_4112; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4114 = 10'h312 == io_inputs_1 ? 7'h0 : _GEN_4113; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4115 = 10'h313 == io_inputs_1 ? 7'h0 : _GEN_4114; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4116 = 10'h314 == io_inputs_1 ? 7'h0 : _GEN_4115; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4117 = 10'h315 == io_inputs_1 ? 7'h0 : _GEN_4116; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4118 = 10'h316 == io_inputs_1 ? 7'h0 : _GEN_4117; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4119 = 10'h317 == io_inputs_1 ? 7'h0 : _GEN_4118; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4120 = 10'h318 == io_inputs_1 ? 7'h0 : _GEN_4119; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4121 = 10'h319 == io_inputs_1 ? 7'h0 : _GEN_4120; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4122 = 10'h31a == io_inputs_1 ? 7'h0 : _GEN_4121; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4123 = 10'h31b == io_inputs_1 ? 7'h0 : _GEN_4122; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4124 = 10'h31c == io_inputs_1 ? 7'h0 : _GEN_4123; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4125 = 10'h31d == io_inputs_1 ? 7'h0 : _GEN_4124; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4126 = 10'h31e == io_inputs_1 ? 7'h0 : _GEN_4125; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4127 = 10'h31f == io_inputs_1 ? 7'h0 : _GEN_4126; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4128 = 10'h320 == io_inputs_1 ? 7'h0 : _GEN_4127; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4129 = 10'h321 == io_inputs_1 ? 7'h0 : _GEN_4128; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4130 = 10'h322 == io_inputs_1 ? 7'h0 : _GEN_4129; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4131 = 10'h323 == io_inputs_1 ? 7'h0 : _GEN_4130; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4132 = 10'h324 == io_inputs_1 ? 7'h0 : _GEN_4131; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4133 = 10'h325 == io_inputs_1 ? 7'h0 : _GEN_4132; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4134 = 10'h326 == io_inputs_1 ? 7'h0 : _GEN_4133; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4135 = 10'h327 == io_inputs_1 ? 7'h0 : _GEN_4134; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4136 = 10'h328 == io_inputs_1 ? 7'h0 : _GEN_4135; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4137 = 10'h329 == io_inputs_1 ? 7'h0 : _GEN_4136; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4138 = 10'h32a == io_inputs_1 ? 7'h0 : _GEN_4137; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4139 = 10'h32b == io_inputs_1 ? 7'h0 : _GEN_4138; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4140 = 10'h32c == io_inputs_1 ? 7'h0 : _GEN_4139; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4141 = 10'h32d == io_inputs_1 ? 7'h0 : _GEN_4140; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4142 = 10'h32e == io_inputs_1 ? 7'h0 : _GEN_4141; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4143 = 10'h32f == io_inputs_1 ? 7'h0 : _GEN_4142; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4144 = 10'h330 == io_inputs_1 ? 7'h0 : _GEN_4143; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4145 = 10'h331 == io_inputs_1 ? 7'h0 : _GEN_4144; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4146 = 10'h332 == io_inputs_1 ? 7'h0 : _GEN_4145; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4147 = 10'h333 == io_inputs_1 ? 7'h0 : _GEN_4146; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4148 = 10'h334 == io_inputs_1 ? 7'h0 : _GEN_4147; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4149 = 10'h335 == io_inputs_1 ? 7'h0 : _GEN_4148; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4150 = 10'h336 == io_inputs_1 ? 7'h0 : _GEN_4149; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4151 = 10'h337 == io_inputs_1 ? 7'h0 : _GEN_4150; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4152 = 10'h338 == io_inputs_1 ? 7'h0 : _GEN_4151; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4153 = 10'h339 == io_inputs_1 ? 7'h0 : _GEN_4152; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4154 = 10'h33a == io_inputs_1 ? 7'h0 : _GEN_4153; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4155 = 10'h33b == io_inputs_1 ? 7'h0 : _GEN_4154; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4156 = 10'h33c == io_inputs_1 ? 7'h0 : _GEN_4155; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4157 = 10'h33d == io_inputs_1 ? 7'h0 : _GEN_4156; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4158 = 10'h33e == io_inputs_1 ? 7'h0 : _GEN_4157; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4159 = 10'h33f == io_inputs_1 ? 7'h0 : _GEN_4158; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4160 = 10'h340 == io_inputs_1 ? 7'h0 : _GEN_4159; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4161 = 10'h341 == io_inputs_1 ? 7'h0 : _GEN_4160; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4162 = 10'h342 == io_inputs_1 ? 7'h0 : _GEN_4161; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4163 = 10'h343 == io_inputs_1 ? 7'h0 : _GEN_4162; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4164 = 10'h344 == io_inputs_1 ? 7'h0 : _GEN_4163; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4165 = 10'h345 == io_inputs_1 ? 7'h0 : _GEN_4164; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4166 = 10'h346 == io_inputs_1 ? 7'h0 : _GEN_4165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4167 = 10'h347 == io_inputs_1 ? 7'h0 : _GEN_4166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4168 = 10'h348 == io_inputs_1 ? 7'h0 : _GEN_4167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4169 = 10'h349 == io_inputs_1 ? 7'h0 : _GEN_4168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4170 = 10'h34a == io_inputs_1 ? 7'h0 : _GEN_4169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4171 = 10'h34b == io_inputs_1 ? 7'h0 : _GEN_4170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4172 = 10'h34c == io_inputs_1 ? 7'h0 : _GEN_4171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4173 = 10'h34d == io_inputs_1 ? 7'h0 : _GEN_4172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4174 = 10'h34e == io_inputs_1 ? 7'h0 : _GEN_4173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4175 = 10'h34f == io_inputs_1 ? 7'h0 : _GEN_4174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4176 = 10'h350 == io_inputs_1 ? 7'h0 : _GEN_4175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4177 = 10'h351 == io_inputs_1 ? 7'h0 : _GEN_4176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4178 = 10'h352 == io_inputs_1 ? 7'h0 : _GEN_4177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4179 = 10'h353 == io_inputs_1 ? 7'h0 : _GEN_4178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4180 = 10'h354 == io_inputs_1 ? 7'h0 : _GEN_4179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4181 = 10'h355 == io_inputs_1 ? 7'h0 : _GEN_4180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4182 = 10'h356 == io_inputs_1 ? 7'h0 : _GEN_4181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4183 = 10'h357 == io_inputs_1 ? 7'h0 : _GEN_4182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4184 = 10'h358 == io_inputs_1 ? 7'h0 : _GEN_4183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4185 = 10'h359 == io_inputs_1 ? 7'h0 : _GEN_4184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4186 = 10'h35a == io_inputs_1 ? 7'h0 : _GEN_4185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4187 = 10'h35b == io_inputs_1 ? 7'h0 : _GEN_4186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4188 = 10'h35c == io_inputs_1 ? 7'h0 : _GEN_4187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4189 = 10'h35d == io_inputs_1 ? 7'h0 : _GEN_4188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4190 = 10'h35e == io_inputs_1 ? 7'h0 : _GEN_4189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4191 = 10'h35f == io_inputs_1 ? 7'h0 : _GEN_4190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4192 = 10'h360 == io_inputs_1 ? 7'h0 : _GEN_4191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4193 = 10'h361 == io_inputs_1 ? 7'h0 : _GEN_4192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4194 = 10'h362 == io_inputs_1 ? 7'h0 : _GEN_4193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4195 = 10'h363 == io_inputs_1 ? 7'h0 : _GEN_4194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4196 = 10'h364 == io_inputs_1 ? 7'h0 : _GEN_4195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4197 = 10'h365 == io_inputs_1 ? 7'h0 : _GEN_4196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4198 = 10'h366 == io_inputs_1 ? 7'h0 : _GEN_4197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4199 = 10'h367 == io_inputs_1 ? 7'h0 : _GEN_4198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4200 = 10'h368 == io_inputs_1 ? 7'h0 : _GEN_4199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4201 = 10'h369 == io_inputs_1 ? 7'h0 : _GEN_4200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4202 = 10'h36a == io_inputs_1 ? 7'h0 : _GEN_4201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4203 = 10'h36b == io_inputs_1 ? 7'h0 : _GEN_4202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4204 = 10'h36c == io_inputs_1 ? 7'h0 : _GEN_4203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4205 = 10'h36d == io_inputs_1 ? 7'h0 : _GEN_4204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4206 = 10'h36e == io_inputs_1 ? 7'h0 : _GEN_4205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4207 = 10'h36f == io_inputs_1 ? 7'h0 : _GEN_4206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4208 = 10'h370 == io_inputs_1 ? 7'h0 : _GEN_4207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4209 = 10'h371 == io_inputs_1 ? 7'h0 : _GEN_4208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4210 = 10'h372 == io_inputs_1 ? 7'h0 : _GEN_4209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4211 = 10'h373 == io_inputs_1 ? 7'h0 : _GEN_4210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4212 = 10'h374 == io_inputs_1 ? 7'h0 : _GEN_4211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4213 = 10'h375 == io_inputs_1 ? 7'h0 : _GEN_4212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4214 = 10'h376 == io_inputs_1 ? 7'h0 : _GEN_4213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4215 = 10'h377 == io_inputs_1 ? 7'h0 : _GEN_4214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4216 = 10'h378 == io_inputs_1 ? 7'h0 : _GEN_4215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4217 = 10'h379 == io_inputs_1 ? 7'h0 : _GEN_4216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4218 = 10'h37a == io_inputs_1 ? 7'h0 : _GEN_4217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4219 = 10'h37b == io_inputs_1 ? 7'h0 : _GEN_4218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4220 = 10'h37c == io_inputs_1 ? 7'h0 : _GEN_4219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4221 = 10'h37d == io_inputs_1 ? 7'h0 : _GEN_4220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4222 = 10'h37e == io_inputs_1 ? 7'h0 : _GEN_4221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4223 = 10'h37f == io_inputs_1 ? 7'h0 : _GEN_4222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4224 = 10'h380 == io_inputs_1 ? 7'h0 : _GEN_4223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4225 = 10'h381 == io_inputs_1 ? 7'h0 : _GEN_4224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4226 = 10'h382 == io_inputs_1 ? 7'h0 : _GEN_4225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4227 = 10'h383 == io_inputs_1 ? 7'h0 : _GEN_4226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4228 = 10'h384 == io_inputs_1 ? 7'h0 : _GEN_4227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4229 = 10'h385 == io_inputs_1 ? 7'h0 : _GEN_4228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4230 = 10'h386 == io_inputs_1 ? 7'h0 : _GEN_4229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4231 = 10'h387 == io_inputs_1 ? 7'h0 : _GEN_4230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4232 = 10'h388 == io_inputs_1 ? 7'h0 : _GEN_4231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4233 = 10'h389 == io_inputs_1 ? 7'h0 : _GEN_4232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4234 = 10'h38a == io_inputs_1 ? 7'h0 : _GEN_4233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4235 = 10'h38b == io_inputs_1 ? 7'h0 : _GEN_4234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4236 = 10'h38c == io_inputs_1 ? 7'h0 : _GEN_4235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4237 = 10'h38d == io_inputs_1 ? 7'h0 : _GEN_4236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4238 = 10'h38e == io_inputs_1 ? 7'h0 : _GEN_4237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4239 = 10'h38f == io_inputs_1 ? 7'h0 : _GEN_4238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4240 = 10'h390 == io_inputs_1 ? 7'h0 : _GEN_4239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4241 = 10'h391 == io_inputs_1 ? 7'h0 : _GEN_4240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4242 = 10'h392 == io_inputs_1 ? 7'h0 : _GEN_4241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4243 = 10'h393 == io_inputs_1 ? 7'h0 : _GEN_4242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4244 = 10'h394 == io_inputs_1 ? 7'h0 : _GEN_4243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4245 = 10'h395 == io_inputs_1 ? 7'h0 : _GEN_4244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4246 = 10'h396 == io_inputs_1 ? 7'h0 : _GEN_4245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4247 = 10'h397 == io_inputs_1 ? 7'h0 : _GEN_4246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4248 = 10'h398 == io_inputs_1 ? 7'h0 : _GEN_4247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4249 = 10'h399 == io_inputs_1 ? 7'h0 : _GEN_4248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4250 = 10'h39a == io_inputs_1 ? 7'h0 : _GEN_4249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4251 = 10'h39b == io_inputs_1 ? 7'h0 : _GEN_4250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4252 = 10'h39c == io_inputs_1 ? 7'h0 : _GEN_4251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4253 = 10'h39d == io_inputs_1 ? 7'h0 : _GEN_4252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4254 = 10'h39e == io_inputs_1 ? 7'h0 : _GEN_4253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4255 = 10'h39f == io_inputs_1 ? 7'h0 : _GEN_4254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4256 = 10'h3a0 == io_inputs_1 ? 7'h0 : _GEN_4255; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4257 = 10'h3a1 == io_inputs_1 ? 7'h0 : _GEN_4256; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4258 = 10'h3a2 == io_inputs_1 ? 7'h0 : _GEN_4257; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4259 = 10'h3a3 == io_inputs_1 ? 7'h0 : _GEN_4258; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4260 = 10'h3a4 == io_inputs_1 ? 7'h0 : _GEN_4259; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4261 = 10'h3a5 == io_inputs_1 ? 7'h0 : _GEN_4260; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4262 = 10'h3a6 == io_inputs_1 ? 7'h0 : _GEN_4261; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4263 = 10'h3a7 == io_inputs_1 ? 7'h0 : _GEN_4262; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4264 = 10'h3a8 == io_inputs_1 ? 7'h0 : _GEN_4263; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4265 = 10'h3a9 == io_inputs_1 ? 7'h0 : _GEN_4264; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4266 = 10'h3aa == io_inputs_1 ? 7'h0 : _GEN_4265; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4267 = 10'h3ab == io_inputs_1 ? 7'h0 : _GEN_4266; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4268 = 10'h3ac == io_inputs_1 ? 7'h0 : _GEN_4267; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4269 = 10'h3ad == io_inputs_1 ? 7'h0 : _GEN_4268; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4270 = 10'h3ae == io_inputs_1 ? 7'h0 : _GEN_4269; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4271 = 10'h3af == io_inputs_1 ? 7'h0 : _GEN_4270; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4272 = 10'h3b0 == io_inputs_1 ? 7'h0 : _GEN_4271; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4273 = 10'h3b1 == io_inputs_1 ? 7'h0 : _GEN_4272; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4274 = 10'h3b2 == io_inputs_1 ? 7'h0 : _GEN_4273; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4275 = 10'h3b3 == io_inputs_1 ? 7'h0 : _GEN_4274; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4276 = 10'h3b4 == io_inputs_1 ? 7'h0 : _GEN_4275; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4277 = 10'h3b5 == io_inputs_1 ? 7'h0 : _GEN_4276; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4278 = 10'h3b6 == io_inputs_1 ? 7'h0 : _GEN_4277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4279 = 10'h3b7 == io_inputs_1 ? 7'h0 : _GEN_4278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4280 = 10'h3b8 == io_inputs_1 ? 7'h0 : _GEN_4279; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4281 = 10'h3b9 == io_inputs_1 ? 7'h0 : _GEN_4280; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4282 = 10'h3ba == io_inputs_1 ? 7'h0 : _GEN_4281; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4283 = 10'h3bb == io_inputs_1 ? 7'h0 : _GEN_4282; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4284 = 10'h3bc == io_inputs_1 ? 7'h0 : _GEN_4283; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4285 = 10'h3bd == io_inputs_1 ? 7'h0 : _GEN_4284; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4286 = 10'h3be == io_inputs_1 ? 7'h0 : _GEN_4285; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4287 = 10'h3bf == io_inputs_1 ? 7'h0 : _GEN_4286; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4288 = 10'h3c0 == io_inputs_1 ? 7'h0 : _GEN_4287; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4289 = 10'h3c1 == io_inputs_1 ? 7'h0 : _GEN_4288; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4290 = 10'h3c2 == io_inputs_1 ? 7'h0 : _GEN_4289; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4291 = 10'h3c3 == io_inputs_1 ? 7'h0 : _GEN_4290; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4292 = 10'h3c4 == io_inputs_1 ? 7'h0 : _GEN_4291; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4293 = 10'h3c5 == io_inputs_1 ? 7'h0 : _GEN_4292; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4294 = 10'h3c6 == io_inputs_1 ? 7'h0 : _GEN_4293; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4295 = 10'h3c7 == io_inputs_1 ? 7'h0 : _GEN_4294; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4296 = 10'h3c8 == io_inputs_1 ? 7'h0 : _GEN_4295; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4297 = 10'h3c9 == io_inputs_1 ? 7'h0 : _GEN_4296; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4298 = 10'h3ca == io_inputs_1 ? 7'h0 : _GEN_4297; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4299 = 10'h3cb == io_inputs_1 ? 7'h0 : _GEN_4298; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4300 = 10'h3cc == io_inputs_1 ? 7'h0 : _GEN_4299; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4301 = 10'h3cd == io_inputs_1 ? 7'h0 : _GEN_4300; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4302 = 10'h3ce == io_inputs_1 ? 7'h0 : _GEN_4301; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4303 = 10'h3cf == io_inputs_1 ? 7'h0 : _GEN_4302; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4304 = 10'h3d0 == io_inputs_1 ? 7'h0 : _GEN_4303; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4305 = 10'h3d1 == io_inputs_1 ? 7'h0 : _GEN_4304; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4306 = 10'h3d2 == io_inputs_1 ? 7'h0 : _GEN_4305; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4307 = 10'h3d3 == io_inputs_1 ? 7'h0 : _GEN_4306; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4308 = 10'h3d4 == io_inputs_1 ? 7'h0 : _GEN_4307; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4309 = 10'h3d5 == io_inputs_1 ? 7'h0 : _GEN_4308; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4310 = 10'h3d6 == io_inputs_1 ? 7'h0 : _GEN_4309; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4311 = 10'h3d7 == io_inputs_1 ? 7'h0 : _GEN_4310; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4312 = 10'h3d8 == io_inputs_1 ? 7'h0 : _GEN_4311; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4313 = 10'h3d9 == io_inputs_1 ? 7'h0 : _GEN_4312; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4314 = 10'h3da == io_inputs_1 ? 7'h0 : _GEN_4313; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4315 = 10'h3db == io_inputs_1 ? 7'h0 : _GEN_4314; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4316 = 10'h3dc == io_inputs_1 ? 7'h0 : _GEN_4315; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4317 = 10'h3dd == io_inputs_1 ? 7'h0 : _GEN_4316; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4318 = 10'h3de == io_inputs_1 ? 7'h0 : _GEN_4317; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4319 = 10'h3df == io_inputs_1 ? 7'h0 : _GEN_4318; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4320 = 10'h3e0 == io_inputs_1 ? 7'h0 : _GEN_4319; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4321 = 10'h3e1 == io_inputs_1 ? 7'h0 : _GEN_4320; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4322 = 10'h3e2 == io_inputs_1 ? 7'h0 : _GEN_4321; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4323 = 10'h3e3 == io_inputs_1 ? 7'h0 : _GEN_4322; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4324 = 10'h3e4 == io_inputs_1 ? 7'h0 : _GEN_4323; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4325 = 10'h3e5 == io_inputs_1 ? 7'h0 : _GEN_4324; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4326 = 10'h3e6 == io_inputs_1 ? 7'h0 : _GEN_4325; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4327 = 10'h3e7 == io_inputs_1 ? 7'h0 : _GEN_4326; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4328 = 10'h3e8 == io_inputs_1 ? 7'h0 : _GEN_4327; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4329 = 10'h3e9 == io_inputs_1 ? 7'h0 : _GEN_4328; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4330 = 10'h3ea == io_inputs_1 ? 7'h0 : _GEN_4329; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4331 = 10'h3eb == io_inputs_1 ? 7'h0 : _GEN_4330; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4332 = 10'h3ec == io_inputs_1 ? 7'h0 : _GEN_4331; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4333 = 10'h3ed == io_inputs_1 ? 7'h0 : _GEN_4332; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4334 = 10'h3ee == io_inputs_1 ? 7'h0 : _GEN_4333; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4335 = 10'h3ef == io_inputs_1 ? 7'h0 : _GEN_4334; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4336 = 10'h3f0 == io_inputs_1 ? 7'h0 : _GEN_4335; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4337 = 10'h3f1 == io_inputs_1 ? 7'h0 : _GEN_4336; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4338 = 10'h3f2 == io_inputs_1 ? 7'h0 : _GEN_4337; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4339 = 10'h3f3 == io_inputs_1 ? 7'h0 : _GEN_4338; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4340 = 10'h3f4 == io_inputs_1 ? 7'h0 : _GEN_4339; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4341 = 10'h3f5 == io_inputs_1 ? 7'h0 : _GEN_4340; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4342 = 10'h3f6 == io_inputs_1 ? 7'h0 : _GEN_4341; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4343 = 10'h3f7 == io_inputs_1 ? 7'h0 : _GEN_4342; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4344 = 10'h3f8 == io_inputs_1 ? 7'h0 : _GEN_4343; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4345 = 10'h3f9 == io_inputs_1 ? 7'h0 : _GEN_4344; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4346 = 10'h3fa == io_inputs_1 ? 7'h0 : _GEN_4345; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4347 = 10'h3fb == io_inputs_1 ? 7'h0 : _GEN_4346; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4348 = 10'h3fc == io_inputs_1 ? 7'h0 : _GEN_4347; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4349 = 10'h3fd == io_inputs_1 ? 7'h0 : _GEN_4348; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4350 = 10'h3fe == io_inputs_1 ? 7'h0 : _GEN_4349; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4351 = 10'h3ff == io_inputs_1 ? 7'h0 : _GEN_4350; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4703 = 10'h15f == io_inputs_1 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4704 = 10'h160 == io_inputs_1 ? 7'h2 : _GEN_4703; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4705 = 10'h161 == io_inputs_1 ? 7'h3 : _GEN_4704; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4706 = 10'h162 == io_inputs_1 ? 7'h4 : _GEN_4705; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4707 = 10'h163 == io_inputs_1 ? 7'h5 : _GEN_4706; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4708 = 10'h164 == io_inputs_1 ? 7'h6 : _GEN_4707; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4709 = 10'h165 == io_inputs_1 ? 7'h7 : _GEN_4708; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4710 = 10'h166 == io_inputs_1 ? 7'h8 : _GEN_4709; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4711 = 10'h167 == io_inputs_1 ? 7'h9 : _GEN_4710; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4712 = 10'h168 == io_inputs_1 ? 7'ha : _GEN_4711; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4713 = 10'h169 == io_inputs_1 ? 7'hb : _GEN_4712; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4714 = 10'h16a == io_inputs_1 ? 7'hc : _GEN_4713; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4715 = 10'h16b == io_inputs_1 ? 7'hd : _GEN_4714; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4716 = 10'h16c == io_inputs_1 ? 7'he : _GEN_4715; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4717 = 10'h16d == io_inputs_1 ? 7'hf : _GEN_4716; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4718 = 10'h16e == io_inputs_1 ? 7'h10 : _GEN_4717; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4719 = 10'h16f == io_inputs_1 ? 7'h11 : _GEN_4718; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4720 = 10'h170 == io_inputs_1 ? 7'h12 : _GEN_4719; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4721 = 10'h171 == io_inputs_1 ? 7'h13 : _GEN_4720; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4722 = 10'h172 == io_inputs_1 ? 7'h14 : _GEN_4721; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4723 = 10'h173 == io_inputs_1 ? 7'h15 : _GEN_4722; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4724 = 10'h174 == io_inputs_1 ? 7'h16 : _GEN_4723; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4725 = 10'h175 == io_inputs_1 ? 7'h17 : _GEN_4724; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4726 = 10'h176 == io_inputs_1 ? 7'h18 : _GEN_4725; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4727 = 10'h177 == io_inputs_1 ? 7'h19 : _GEN_4726; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4728 = 10'h178 == io_inputs_1 ? 7'h1a : _GEN_4727; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4729 = 10'h179 == io_inputs_1 ? 7'h1b : _GEN_4728; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4730 = 10'h17a == io_inputs_1 ? 7'h1c : _GEN_4729; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4731 = 10'h17b == io_inputs_1 ? 7'h1d : _GEN_4730; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4732 = 10'h17c == io_inputs_1 ? 7'h1e : _GEN_4731; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4733 = 10'h17d == io_inputs_1 ? 7'h1f : _GEN_4732; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4734 = 10'h17e == io_inputs_1 ? 7'h20 : _GEN_4733; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4735 = 10'h17f == io_inputs_1 ? 7'h21 : _GEN_4734; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4736 = 10'h180 == io_inputs_1 ? 7'h22 : _GEN_4735; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4737 = 10'h181 == io_inputs_1 ? 7'h23 : _GEN_4736; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4738 = 10'h182 == io_inputs_1 ? 7'h24 : _GEN_4737; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4739 = 10'h183 == io_inputs_1 ? 7'h25 : _GEN_4738; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4740 = 10'h184 == io_inputs_1 ? 7'h26 : _GEN_4739; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4741 = 10'h185 == io_inputs_1 ? 7'h27 : _GEN_4740; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4742 = 10'h186 == io_inputs_1 ? 7'h28 : _GEN_4741; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4743 = 10'h187 == io_inputs_1 ? 7'h29 : _GEN_4742; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4744 = 10'h188 == io_inputs_1 ? 7'h2a : _GEN_4743; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4745 = 10'h189 == io_inputs_1 ? 7'h2b : _GEN_4744; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4746 = 10'h18a == io_inputs_1 ? 7'h2c : _GEN_4745; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4747 = 10'h18b == io_inputs_1 ? 7'h2d : _GEN_4746; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4748 = 10'h18c == io_inputs_1 ? 7'h2e : _GEN_4747; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4749 = 10'h18d == io_inputs_1 ? 7'h2f : _GEN_4748; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4750 = 10'h18e == io_inputs_1 ? 7'h30 : _GEN_4749; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4751 = 10'h18f == io_inputs_1 ? 7'h31 : _GEN_4750; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4752 = 10'h190 == io_inputs_1 ? 7'h32 : _GEN_4751; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4753 = 10'h191 == io_inputs_1 ? 7'h33 : _GEN_4752; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4754 = 10'h192 == io_inputs_1 ? 7'h34 : _GEN_4753; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4755 = 10'h193 == io_inputs_1 ? 7'h35 : _GEN_4754; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4756 = 10'h194 == io_inputs_1 ? 7'h36 : _GEN_4755; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4757 = 10'h195 == io_inputs_1 ? 7'h37 : _GEN_4756; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4758 = 10'h196 == io_inputs_1 ? 7'h38 : _GEN_4757; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4759 = 10'h197 == io_inputs_1 ? 7'h39 : _GEN_4758; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4760 = 10'h198 == io_inputs_1 ? 7'h3a : _GEN_4759; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4761 = 10'h199 == io_inputs_1 ? 7'h3b : _GEN_4760; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4762 = 10'h19a == io_inputs_1 ? 7'h3c : _GEN_4761; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4763 = 10'h19b == io_inputs_1 ? 7'h3d : _GEN_4762; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4764 = 10'h19c == io_inputs_1 ? 7'h3e : _GEN_4763; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4765 = 10'h19d == io_inputs_1 ? 7'h3f : _GEN_4764; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4766 = 10'h19e == io_inputs_1 ? 7'h40 : _GEN_4765; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4767 = 10'h19f == io_inputs_1 ? 7'h41 : _GEN_4766; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4768 = 10'h1a0 == io_inputs_1 ? 7'h42 : _GEN_4767; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4769 = 10'h1a1 == io_inputs_1 ? 7'h43 : _GEN_4768; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4770 = 10'h1a2 == io_inputs_1 ? 7'h44 : _GEN_4769; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4771 = 10'h1a3 == io_inputs_1 ? 7'h45 : _GEN_4770; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4772 = 10'h1a4 == io_inputs_1 ? 7'h46 : _GEN_4771; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4773 = 10'h1a5 == io_inputs_1 ? 7'h47 : _GEN_4772; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4774 = 10'h1a6 == io_inputs_1 ? 7'h48 : _GEN_4773; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4775 = 10'h1a7 == io_inputs_1 ? 7'h49 : _GEN_4774; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4776 = 10'h1a8 == io_inputs_1 ? 7'h4a : _GEN_4775; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4777 = 10'h1a9 == io_inputs_1 ? 7'h4b : _GEN_4776; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4778 = 10'h1aa == io_inputs_1 ? 7'h4c : _GEN_4777; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4779 = 10'h1ab == io_inputs_1 ? 7'h4d : _GEN_4778; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4780 = 10'h1ac == io_inputs_1 ? 7'h4e : _GEN_4779; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4781 = 10'h1ad == io_inputs_1 ? 7'h4f : _GEN_4780; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4782 = 10'h1ae == io_inputs_1 ? 7'h50 : _GEN_4781; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4783 = 10'h1af == io_inputs_1 ? 7'h51 : _GEN_4782; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4784 = 10'h1b0 == io_inputs_1 ? 7'h52 : _GEN_4783; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4785 = 10'h1b1 == io_inputs_1 ? 7'h53 : _GEN_4784; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4786 = 10'h1b2 == io_inputs_1 ? 7'h54 : _GEN_4785; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4787 = 10'h1b3 == io_inputs_1 ? 7'h55 : _GEN_4786; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4788 = 10'h1b4 == io_inputs_1 ? 7'h56 : _GEN_4787; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4789 = 10'h1b5 == io_inputs_1 ? 7'h57 : _GEN_4788; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4790 = 10'h1b6 == io_inputs_1 ? 7'h58 : _GEN_4789; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4791 = 10'h1b7 == io_inputs_1 ? 7'h59 : _GEN_4790; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4792 = 10'h1b8 == io_inputs_1 ? 7'h5a : _GEN_4791; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4793 = 10'h1b9 == io_inputs_1 ? 7'h5b : _GEN_4792; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4794 = 10'h1ba == io_inputs_1 ? 7'h5c : _GEN_4793; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4795 = 10'h1bb == io_inputs_1 ? 7'h5d : _GEN_4794; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4796 = 10'h1bc == io_inputs_1 ? 7'h5e : _GEN_4795; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4797 = 10'h1bd == io_inputs_1 ? 7'h5f : _GEN_4796; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4798 = 10'h1be == io_inputs_1 ? 7'h60 : _GEN_4797; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4799 = 10'h1bf == io_inputs_1 ? 7'h61 : _GEN_4798; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4800 = 10'h1c0 == io_inputs_1 ? 7'h62 : _GEN_4799; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4801 = 10'h1c1 == io_inputs_1 ? 7'h63 : _GEN_4800; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4802 = 10'h1c2 == io_inputs_1 ? 7'h64 : _GEN_4801; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4803 = 10'h1c3 == io_inputs_1 ? 7'h63 : _GEN_4802; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4804 = 10'h1c4 == io_inputs_1 ? 7'h62 : _GEN_4803; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4805 = 10'h1c5 == io_inputs_1 ? 7'h61 : _GEN_4804; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4806 = 10'h1c6 == io_inputs_1 ? 7'h60 : _GEN_4805; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4807 = 10'h1c7 == io_inputs_1 ? 7'h5f : _GEN_4806; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4808 = 10'h1c8 == io_inputs_1 ? 7'h5e : _GEN_4807; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4809 = 10'h1c9 == io_inputs_1 ? 7'h5d : _GEN_4808; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4810 = 10'h1ca == io_inputs_1 ? 7'h5c : _GEN_4809; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4811 = 10'h1cb == io_inputs_1 ? 7'h5b : _GEN_4810; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4812 = 10'h1cc == io_inputs_1 ? 7'h5a : _GEN_4811; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4813 = 10'h1cd == io_inputs_1 ? 7'h59 : _GEN_4812; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4814 = 10'h1ce == io_inputs_1 ? 7'h58 : _GEN_4813; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4815 = 10'h1cf == io_inputs_1 ? 7'h57 : _GEN_4814; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4816 = 10'h1d0 == io_inputs_1 ? 7'h56 : _GEN_4815; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4817 = 10'h1d1 == io_inputs_1 ? 7'h55 : _GEN_4816; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4818 = 10'h1d2 == io_inputs_1 ? 7'h54 : _GEN_4817; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4819 = 10'h1d3 == io_inputs_1 ? 7'h53 : _GEN_4818; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4820 = 10'h1d4 == io_inputs_1 ? 7'h52 : _GEN_4819; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4821 = 10'h1d5 == io_inputs_1 ? 7'h51 : _GEN_4820; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4822 = 10'h1d6 == io_inputs_1 ? 7'h50 : _GEN_4821; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4823 = 10'h1d7 == io_inputs_1 ? 7'h4f : _GEN_4822; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4824 = 10'h1d8 == io_inputs_1 ? 7'h4e : _GEN_4823; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4825 = 10'h1d9 == io_inputs_1 ? 7'h4d : _GEN_4824; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4826 = 10'h1da == io_inputs_1 ? 7'h4c : _GEN_4825; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4827 = 10'h1db == io_inputs_1 ? 7'h4b : _GEN_4826; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4828 = 10'h1dc == io_inputs_1 ? 7'h4a : _GEN_4827; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4829 = 10'h1dd == io_inputs_1 ? 7'h49 : _GEN_4828; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4830 = 10'h1de == io_inputs_1 ? 7'h48 : _GEN_4829; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4831 = 10'h1df == io_inputs_1 ? 7'h47 : _GEN_4830; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4832 = 10'h1e0 == io_inputs_1 ? 7'h46 : _GEN_4831; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4833 = 10'h1e1 == io_inputs_1 ? 7'h45 : _GEN_4832; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4834 = 10'h1e2 == io_inputs_1 ? 7'h44 : _GEN_4833; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4835 = 10'h1e3 == io_inputs_1 ? 7'h43 : _GEN_4834; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4836 = 10'h1e4 == io_inputs_1 ? 7'h42 : _GEN_4835; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4837 = 10'h1e5 == io_inputs_1 ? 7'h41 : _GEN_4836; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4838 = 10'h1e6 == io_inputs_1 ? 7'h40 : _GEN_4837; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4839 = 10'h1e7 == io_inputs_1 ? 7'h3f : _GEN_4838; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4840 = 10'h1e8 == io_inputs_1 ? 7'h3e : _GEN_4839; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4841 = 10'h1e9 == io_inputs_1 ? 7'h3d : _GEN_4840; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4842 = 10'h1ea == io_inputs_1 ? 7'h3c : _GEN_4841; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4843 = 10'h1eb == io_inputs_1 ? 7'h3b : _GEN_4842; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4844 = 10'h1ec == io_inputs_1 ? 7'h3a : _GEN_4843; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4845 = 10'h1ed == io_inputs_1 ? 7'h39 : _GEN_4844; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4846 = 10'h1ee == io_inputs_1 ? 7'h38 : _GEN_4845; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4847 = 10'h1ef == io_inputs_1 ? 7'h37 : _GEN_4846; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4848 = 10'h1f0 == io_inputs_1 ? 7'h36 : _GEN_4847; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4849 = 10'h1f1 == io_inputs_1 ? 7'h35 : _GEN_4848; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4850 = 10'h1f2 == io_inputs_1 ? 7'h34 : _GEN_4849; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4851 = 10'h1f3 == io_inputs_1 ? 7'h33 : _GEN_4850; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4852 = 10'h1f4 == io_inputs_1 ? 7'h32 : _GEN_4851; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4853 = 10'h1f5 == io_inputs_1 ? 7'h31 : _GEN_4852; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4854 = 10'h1f6 == io_inputs_1 ? 7'h30 : _GEN_4853; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4855 = 10'h1f7 == io_inputs_1 ? 7'h2f : _GEN_4854; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4856 = 10'h1f8 == io_inputs_1 ? 7'h2e : _GEN_4855; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4857 = 10'h1f9 == io_inputs_1 ? 7'h2d : _GEN_4856; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4858 = 10'h1fa == io_inputs_1 ? 7'h2c : _GEN_4857; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4859 = 10'h1fb == io_inputs_1 ? 7'h2b : _GEN_4858; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4860 = 10'h1fc == io_inputs_1 ? 7'h2a : _GEN_4859; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4861 = 10'h1fd == io_inputs_1 ? 7'h29 : _GEN_4860; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4862 = 10'h1fe == io_inputs_1 ? 7'h28 : _GEN_4861; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4863 = 10'h1ff == io_inputs_1 ? 7'h27 : _GEN_4862; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4864 = 10'h200 == io_inputs_1 ? 7'h26 : _GEN_4863; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4865 = 10'h201 == io_inputs_1 ? 7'h25 : _GEN_4864; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4866 = 10'h202 == io_inputs_1 ? 7'h24 : _GEN_4865; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4867 = 10'h203 == io_inputs_1 ? 7'h23 : _GEN_4866; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4868 = 10'h204 == io_inputs_1 ? 7'h22 : _GEN_4867; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4869 = 10'h205 == io_inputs_1 ? 7'h21 : _GEN_4868; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4870 = 10'h206 == io_inputs_1 ? 7'h20 : _GEN_4869; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4871 = 10'h207 == io_inputs_1 ? 7'h1f : _GEN_4870; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4872 = 10'h208 == io_inputs_1 ? 7'h1e : _GEN_4871; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4873 = 10'h209 == io_inputs_1 ? 7'h1d : _GEN_4872; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4874 = 10'h20a == io_inputs_1 ? 7'h1c : _GEN_4873; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4875 = 10'h20b == io_inputs_1 ? 7'h1b : _GEN_4874; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4876 = 10'h20c == io_inputs_1 ? 7'h1a : _GEN_4875; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4877 = 10'h20d == io_inputs_1 ? 7'h19 : _GEN_4876; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4878 = 10'h20e == io_inputs_1 ? 7'h18 : _GEN_4877; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4879 = 10'h20f == io_inputs_1 ? 7'h17 : _GEN_4878; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4880 = 10'h210 == io_inputs_1 ? 7'h16 : _GEN_4879; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4881 = 10'h211 == io_inputs_1 ? 7'h15 : _GEN_4880; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4882 = 10'h212 == io_inputs_1 ? 7'h14 : _GEN_4881; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4883 = 10'h213 == io_inputs_1 ? 7'h13 : _GEN_4882; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4884 = 10'h214 == io_inputs_1 ? 7'h12 : _GEN_4883; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4885 = 10'h215 == io_inputs_1 ? 7'h11 : _GEN_4884; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4886 = 10'h216 == io_inputs_1 ? 7'h10 : _GEN_4885; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4887 = 10'h217 == io_inputs_1 ? 7'hf : _GEN_4886; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4888 = 10'h218 == io_inputs_1 ? 7'he : _GEN_4887; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4889 = 10'h219 == io_inputs_1 ? 7'hd : _GEN_4888; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4890 = 10'h21a == io_inputs_1 ? 7'hc : _GEN_4889; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4891 = 10'h21b == io_inputs_1 ? 7'hb : _GEN_4890; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4892 = 10'h21c == io_inputs_1 ? 7'ha : _GEN_4891; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4893 = 10'h21d == io_inputs_1 ? 7'h9 : _GEN_4892; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4894 = 10'h21e == io_inputs_1 ? 7'h8 : _GEN_4893; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4895 = 10'h21f == io_inputs_1 ? 7'h7 : _GEN_4894; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4896 = 10'h220 == io_inputs_1 ? 7'h6 : _GEN_4895; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4897 = 10'h221 == io_inputs_1 ? 7'h5 : _GEN_4896; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4898 = 10'h222 == io_inputs_1 ? 7'h4 : _GEN_4897; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4899 = 10'h223 == io_inputs_1 ? 7'h3 : _GEN_4898; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4900 = 10'h224 == io_inputs_1 ? 7'h2 : _GEN_4899; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4901 = 10'h225 == io_inputs_1 ? 7'h1 : _GEN_4900; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4902 = 10'h226 == io_inputs_1 ? 7'h0 : _GEN_4901; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4903 = 10'h227 == io_inputs_1 ? 7'h0 : _GEN_4902; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4904 = 10'h228 == io_inputs_1 ? 7'h0 : _GEN_4903; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4905 = 10'h229 == io_inputs_1 ? 7'h0 : _GEN_4904; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4906 = 10'h22a == io_inputs_1 ? 7'h0 : _GEN_4905; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4907 = 10'h22b == io_inputs_1 ? 7'h0 : _GEN_4906; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4908 = 10'h22c == io_inputs_1 ? 7'h0 : _GEN_4907; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4909 = 10'h22d == io_inputs_1 ? 7'h0 : _GEN_4908; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4910 = 10'h22e == io_inputs_1 ? 7'h0 : _GEN_4909; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4911 = 10'h22f == io_inputs_1 ? 7'h0 : _GEN_4910; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4912 = 10'h230 == io_inputs_1 ? 7'h0 : _GEN_4911; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4913 = 10'h231 == io_inputs_1 ? 7'h0 : _GEN_4912; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4914 = 10'h232 == io_inputs_1 ? 7'h0 : _GEN_4913; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4915 = 10'h233 == io_inputs_1 ? 7'h0 : _GEN_4914; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4916 = 10'h234 == io_inputs_1 ? 7'h0 : _GEN_4915; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4917 = 10'h235 == io_inputs_1 ? 7'h0 : _GEN_4916; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4918 = 10'h236 == io_inputs_1 ? 7'h0 : _GEN_4917; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4919 = 10'h237 == io_inputs_1 ? 7'h0 : _GEN_4918; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4920 = 10'h238 == io_inputs_1 ? 7'h0 : _GEN_4919; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4921 = 10'h239 == io_inputs_1 ? 7'h0 : _GEN_4920; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4922 = 10'h23a == io_inputs_1 ? 7'h0 : _GEN_4921; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4923 = 10'h23b == io_inputs_1 ? 7'h0 : _GEN_4922; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4924 = 10'h23c == io_inputs_1 ? 7'h0 : _GEN_4923; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4925 = 10'h23d == io_inputs_1 ? 7'h0 : _GEN_4924; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4926 = 10'h23e == io_inputs_1 ? 7'h0 : _GEN_4925; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4927 = 10'h23f == io_inputs_1 ? 7'h0 : _GEN_4926; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4928 = 10'h240 == io_inputs_1 ? 7'h0 : _GEN_4927; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4929 = 10'h241 == io_inputs_1 ? 7'h0 : _GEN_4928; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4930 = 10'h242 == io_inputs_1 ? 7'h0 : _GEN_4929; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4931 = 10'h243 == io_inputs_1 ? 7'h0 : _GEN_4930; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4932 = 10'h244 == io_inputs_1 ? 7'h0 : _GEN_4931; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4933 = 10'h245 == io_inputs_1 ? 7'h0 : _GEN_4932; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4934 = 10'h246 == io_inputs_1 ? 7'h0 : _GEN_4933; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4935 = 10'h247 == io_inputs_1 ? 7'h0 : _GEN_4934; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4936 = 10'h248 == io_inputs_1 ? 7'h0 : _GEN_4935; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4937 = 10'h249 == io_inputs_1 ? 7'h0 : _GEN_4936; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4938 = 10'h24a == io_inputs_1 ? 7'h0 : _GEN_4937; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4939 = 10'h24b == io_inputs_1 ? 7'h0 : _GEN_4938; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4940 = 10'h24c == io_inputs_1 ? 7'h0 : _GEN_4939; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4941 = 10'h24d == io_inputs_1 ? 7'h0 : _GEN_4940; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4942 = 10'h24e == io_inputs_1 ? 7'h0 : _GEN_4941; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4943 = 10'h24f == io_inputs_1 ? 7'h0 : _GEN_4942; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4944 = 10'h250 == io_inputs_1 ? 7'h0 : _GEN_4943; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4945 = 10'h251 == io_inputs_1 ? 7'h0 : _GEN_4944; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4946 = 10'h252 == io_inputs_1 ? 7'h0 : _GEN_4945; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4947 = 10'h253 == io_inputs_1 ? 7'h0 : _GEN_4946; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4948 = 10'h254 == io_inputs_1 ? 7'h0 : _GEN_4947; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4949 = 10'h255 == io_inputs_1 ? 7'h0 : _GEN_4948; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4950 = 10'h256 == io_inputs_1 ? 7'h0 : _GEN_4949; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4951 = 10'h257 == io_inputs_1 ? 7'h0 : _GEN_4950; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4952 = 10'h258 == io_inputs_1 ? 7'h0 : _GEN_4951; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4953 = 10'h259 == io_inputs_1 ? 7'h0 : _GEN_4952; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4954 = 10'h25a == io_inputs_1 ? 7'h0 : _GEN_4953; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4955 = 10'h25b == io_inputs_1 ? 7'h0 : _GEN_4954; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4956 = 10'h25c == io_inputs_1 ? 7'h0 : _GEN_4955; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4957 = 10'h25d == io_inputs_1 ? 7'h0 : _GEN_4956; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4958 = 10'h25e == io_inputs_1 ? 7'h0 : _GEN_4957; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4959 = 10'h25f == io_inputs_1 ? 7'h0 : _GEN_4958; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4960 = 10'h260 == io_inputs_1 ? 7'h0 : _GEN_4959; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4961 = 10'h261 == io_inputs_1 ? 7'h0 : _GEN_4960; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4962 = 10'h262 == io_inputs_1 ? 7'h0 : _GEN_4961; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4963 = 10'h263 == io_inputs_1 ? 7'h0 : _GEN_4962; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4964 = 10'h264 == io_inputs_1 ? 7'h0 : _GEN_4963; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4965 = 10'h265 == io_inputs_1 ? 7'h0 : _GEN_4964; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4966 = 10'h266 == io_inputs_1 ? 7'h0 : _GEN_4965; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4967 = 10'h267 == io_inputs_1 ? 7'h0 : _GEN_4966; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4968 = 10'h268 == io_inputs_1 ? 7'h0 : _GEN_4967; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4969 = 10'h269 == io_inputs_1 ? 7'h0 : _GEN_4968; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4970 = 10'h26a == io_inputs_1 ? 7'h0 : _GEN_4969; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4971 = 10'h26b == io_inputs_1 ? 7'h0 : _GEN_4970; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4972 = 10'h26c == io_inputs_1 ? 7'h0 : _GEN_4971; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4973 = 10'h26d == io_inputs_1 ? 7'h0 : _GEN_4972; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4974 = 10'h26e == io_inputs_1 ? 7'h0 : _GEN_4973; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4975 = 10'h26f == io_inputs_1 ? 7'h0 : _GEN_4974; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4976 = 10'h270 == io_inputs_1 ? 7'h0 : _GEN_4975; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4977 = 10'h271 == io_inputs_1 ? 7'h0 : _GEN_4976; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4978 = 10'h272 == io_inputs_1 ? 7'h0 : _GEN_4977; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4979 = 10'h273 == io_inputs_1 ? 7'h0 : _GEN_4978; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4980 = 10'h274 == io_inputs_1 ? 7'h0 : _GEN_4979; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4981 = 10'h275 == io_inputs_1 ? 7'h0 : _GEN_4980; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4982 = 10'h276 == io_inputs_1 ? 7'h0 : _GEN_4981; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4983 = 10'h277 == io_inputs_1 ? 7'h0 : _GEN_4982; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4984 = 10'h278 == io_inputs_1 ? 7'h0 : _GEN_4983; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4985 = 10'h279 == io_inputs_1 ? 7'h0 : _GEN_4984; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4986 = 10'h27a == io_inputs_1 ? 7'h0 : _GEN_4985; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4987 = 10'h27b == io_inputs_1 ? 7'h0 : _GEN_4986; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4988 = 10'h27c == io_inputs_1 ? 7'h0 : _GEN_4987; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4989 = 10'h27d == io_inputs_1 ? 7'h0 : _GEN_4988; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4990 = 10'h27e == io_inputs_1 ? 7'h0 : _GEN_4989; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4991 = 10'h27f == io_inputs_1 ? 7'h0 : _GEN_4990; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4992 = 10'h280 == io_inputs_1 ? 7'h0 : _GEN_4991; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4993 = 10'h281 == io_inputs_1 ? 7'h0 : _GEN_4992; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4994 = 10'h282 == io_inputs_1 ? 7'h0 : _GEN_4993; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4995 = 10'h283 == io_inputs_1 ? 7'h0 : _GEN_4994; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4996 = 10'h284 == io_inputs_1 ? 7'h0 : _GEN_4995; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4997 = 10'h285 == io_inputs_1 ? 7'h0 : _GEN_4996; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4998 = 10'h286 == io_inputs_1 ? 7'h0 : _GEN_4997; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_4999 = 10'h287 == io_inputs_1 ? 7'h0 : _GEN_4998; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5000 = 10'h288 == io_inputs_1 ? 7'h0 : _GEN_4999; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5001 = 10'h289 == io_inputs_1 ? 7'h0 : _GEN_5000; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5002 = 10'h28a == io_inputs_1 ? 7'h0 : _GEN_5001; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5003 = 10'h28b == io_inputs_1 ? 7'h0 : _GEN_5002; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5004 = 10'h28c == io_inputs_1 ? 7'h0 : _GEN_5003; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5005 = 10'h28d == io_inputs_1 ? 7'h0 : _GEN_5004; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5006 = 10'h28e == io_inputs_1 ? 7'h0 : _GEN_5005; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5007 = 10'h28f == io_inputs_1 ? 7'h0 : _GEN_5006; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5008 = 10'h290 == io_inputs_1 ? 7'h0 : _GEN_5007; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5009 = 10'h291 == io_inputs_1 ? 7'h0 : _GEN_5008; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5010 = 10'h292 == io_inputs_1 ? 7'h0 : _GEN_5009; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5011 = 10'h293 == io_inputs_1 ? 7'h0 : _GEN_5010; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5012 = 10'h294 == io_inputs_1 ? 7'h0 : _GEN_5011; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5013 = 10'h295 == io_inputs_1 ? 7'h0 : _GEN_5012; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5014 = 10'h296 == io_inputs_1 ? 7'h0 : _GEN_5013; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5015 = 10'h297 == io_inputs_1 ? 7'h0 : _GEN_5014; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5016 = 10'h298 == io_inputs_1 ? 7'h0 : _GEN_5015; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5017 = 10'h299 == io_inputs_1 ? 7'h0 : _GEN_5016; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5018 = 10'h29a == io_inputs_1 ? 7'h0 : _GEN_5017; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5019 = 10'h29b == io_inputs_1 ? 7'h0 : _GEN_5018; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5020 = 10'h29c == io_inputs_1 ? 7'h0 : _GEN_5019; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5021 = 10'h29d == io_inputs_1 ? 7'h0 : _GEN_5020; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5022 = 10'h29e == io_inputs_1 ? 7'h0 : _GEN_5021; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5023 = 10'h29f == io_inputs_1 ? 7'h0 : _GEN_5022; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5024 = 10'h2a0 == io_inputs_1 ? 7'h0 : _GEN_5023; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5025 = 10'h2a1 == io_inputs_1 ? 7'h0 : _GEN_5024; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5026 = 10'h2a2 == io_inputs_1 ? 7'h0 : _GEN_5025; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5027 = 10'h2a3 == io_inputs_1 ? 7'h0 : _GEN_5026; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5028 = 10'h2a4 == io_inputs_1 ? 7'h0 : _GEN_5027; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5029 = 10'h2a5 == io_inputs_1 ? 7'h0 : _GEN_5028; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5030 = 10'h2a6 == io_inputs_1 ? 7'h0 : _GEN_5029; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5031 = 10'h2a7 == io_inputs_1 ? 7'h0 : _GEN_5030; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5032 = 10'h2a8 == io_inputs_1 ? 7'h0 : _GEN_5031; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5033 = 10'h2a9 == io_inputs_1 ? 7'h0 : _GEN_5032; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5034 = 10'h2aa == io_inputs_1 ? 7'h0 : _GEN_5033; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5035 = 10'h2ab == io_inputs_1 ? 7'h0 : _GEN_5034; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5036 = 10'h2ac == io_inputs_1 ? 7'h0 : _GEN_5035; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5037 = 10'h2ad == io_inputs_1 ? 7'h0 : _GEN_5036; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5038 = 10'h2ae == io_inputs_1 ? 7'h0 : _GEN_5037; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5039 = 10'h2af == io_inputs_1 ? 7'h0 : _GEN_5038; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5040 = 10'h2b0 == io_inputs_1 ? 7'h0 : _GEN_5039; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5041 = 10'h2b1 == io_inputs_1 ? 7'h0 : _GEN_5040; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5042 = 10'h2b2 == io_inputs_1 ? 7'h0 : _GEN_5041; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5043 = 10'h2b3 == io_inputs_1 ? 7'h0 : _GEN_5042; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5044 = 10'h2b4 == io_inputs_1 ? 7'h0 : _GEN_5043; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5045 = 10'h2b5 == io_inputs_1 ? 7'h0 : _GEN_5044; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5046 = 10'h2b6 == io_inputs_1 ? 7'h0 : _GEN_5045; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5047 = 10'h2b7 == io_inputs_1 ? 7'h0 : _GEN_5046; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5048 = 10'h2b8 == io_inputs_1 ? 7'h0 : _GEN_5047; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5049 = 10'h2b9 == io_inputs_1 ? 7'h0 : _GEN_5048; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5050 = 10'h2ba == io_inputs_1 ? 7'h0 : _GEN_5049; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5051 = 10'h2bb == io_inputs_1 ? 7'h0 : _GEN_5050; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5052 = 10'h2bc == io_inputs_1 ? 7'h0 : _GEN_5051; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5053 = 10'h2bd == io_inputs_1 ? 7'h0 : _GEN_5052; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5054 = 10'h2be == io_inputs_1 ? 7'h0 : _GEN_5053; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5055 = 10'h2bf == io_inputs_1 ? 7'h0 : _GEN_5054; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5056 = 10'h2c0 == io_inputs_1 ? 7'h0 : _GEN_5055; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5057 = 10'h2c1 == io_inputs_1 ? 7'h0 : _GEN_5056; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5058 = 10'h2c2 == io_inputs_1 ? 7'h0 : _GEN_5057; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5059 = 10'h2c3 == io_inputs_1 ? 7'h0 : _GEN_5058; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5060 = 10'h2c4 == io_inputs_1 ? 7'h0 : _GEN_5059; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5061 = 10'h2c5 == io_inputs_1 ? 7'h0 : _GEN_5060; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5062 = 10'h2c6 == io_inputs_1 ? 7'h0 : _GEN_5061; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5063 = 10'h2c7 == io_inputs_1 ? 7'h0 : _GEN_5062; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5064 = 10'h2c8 == io_inputs_1 ? 7'h0 : _GEN_5063; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5065 = 10'h2c9 == io_inputs_1 ? 7'h0 : _GEN_5064; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5066 = 10'h2ca == io_inputs_1 ? 7'h0 : _GEN_5065; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5067 = 10'h2cb == io_inputs_1 ? 7'h0 : _GEN_5066; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5068 = 10'h2cc == io_inputs_1 ? 7'h0 : _GEN_5067; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5069 = 10'h2cd == io_inputs_1 ? 7'h0 : _GEN_5068; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5070 = 10'h2ce == io_inputs_1 ? 7'h0 : _GEN_5069; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5071 = 10'h2cf == io_inputs_1 ? 7'h0 : _GEN_5070; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5072 = 10'h2d0 == io_inputs_1 ? 7'h0 : _GEN_5071; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5073 = 10'h2d1 == io_inputs_1 ? 7'h0 : _GEN_5072; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5074 = 10'h2d2 == io_inputs_1 ? 7'h0 : _GEN_5073; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5075 = 10'h2d3 == io_inputs_1 ? 7'h0 : _GEN_5074; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5076 = 10'h2d4 == io_inputs_1 ? 7'h0 : _GEN_5075; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5077 = 10'h2d5 == io_inputs_1 ? 7'h0 : _GEN_5076; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5078 = 10'h2d6 == io_inputs_1 ? 7'h0 : _GEN_5077; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5079 = 10'h2d7 == io_inputs_1 ? 7'h0 : _GEN_5078; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5080 = 10'h2d8 == io_inputs_1 ? 7'h0 : _GEN_5079; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5081 = 10'h2d9 == io_inputs_1 ? 7'h0 : _GEN_5080; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5082 = 10'h2da == io_inputs_1 ? 7'h0 : _GEN_5081; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5083 = 10'h2db == io_inputs_1 ? 7'h0 : _GEN_5082; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5084 = 10'h2dc == io_inputs_1 ? 7'h0 : _GEN_5083; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5085 = 10'h2dd == io_inputs_1 ? 7'h0 : _GEN_5084; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5086 = 10'h2de == io_inputs_1 ? 7'h0 : _GEN_5085; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5087 = 10'h2df == io_inputs_1 ? 7'h0 : _GEN_5086; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5088 = 10'h2e0 == io_inputs_1 ? 7'h0 : _GEN_5087; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5089 = 10'h2e1 == io_inputs_1 ? 7'h0 : _GEN_5088; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5090 = 10'h2e2 == io_inputs_1 ? 7'h0 : _GEN_5089; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5091 = 10'h2e3 == io_inputs_1 ? 7'h0 : _GEN_5090; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5092 = 10'h2e4 == io_inputs_1 ? 7'h0 : _GEN_5091; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5093 = 10'h2e5 == io_inputs_1 ? 7'h0 : _GEN_5092; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5094 = 10'h2e6 == io_inputs_1 ? 7'h0 : _GEN_5093; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5095 = 10'h2e7 == io_inputs_1 ? 7'h0 : _GEN_5094; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5096 = 10'h2e8 == io_inputs_1 ? 7'h0 : _GEN_5095; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5097 = 10'h2e9 == io_inputs_1 ? 7'h0 : _GEN_5096; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5098 = 10'h2ea == io_inputs_1 ? 7'h0 : _GEN_5097; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5099 = 10'h2eb == io_inputs_1 ? 7'h0 : _GEN_5098; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5100 = 10'h2ec == io_inputs_1 ? 7'h0 : _GEN_5099; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5101 = 10'h2ed == io_inputs_1 ? 7'h0 : _GEN_5100; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5102 = 10'h2ee == io_inputs_1 ? 7'h0 : _GEN_5101; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5103 = 10'h2ef == io_inputs_1 ? 7'h0 : _GEN_5102; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5104 = 10'h2f0 == io_inputs_1 ? 7'h0 : _GEN_5103; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5105 = 10'h2f1 == io_inputs_1 ? 7'h0 : _GEN_5104; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5106 = 10'h2f2 == io_inputs_1 ? 7'h0 : _GEN_5105; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5107 = 10'h2f3 == io_inputs_1 ? 7'h0 : _GEN_5106; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5108 = 10'h2f4 == io_inputs_1 ? 7'h0 : _GEN_5107; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5109 = 10'h2f5 == io_inputs_1 ? 7'h0 : _GEN_5108; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5110 = 10'h2f6 == io_inputs_1 ? 7'h0 : _GEN_5109; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5111 = 10'h2f7 == io_inputs_1 ? 7'h0 : _GEN_5110; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5112 = 10'h2f8 == io_inputs_1 ? 7'h0 : _GEN_5111; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5113 = 10'h2f9 == io_inputs_1 ? 7'h0 : _GEN_5112; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5114 = 10'h2fa == io_inputs_1 ? 7'h0 : _GEN_5113; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5115 = 10'h2fb == io_inputs_1 ? 7'h0 : _GEN_5114; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5116 = 10'h2fc == io_inputs_1 ? 7'h0 : _GEN_5115; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5117 = 10'h2fd == io_inputs_1 ? 7'h0 : _GEN_5116; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5118 = 10'h2fe == io_inputs_1 ? 7'h0 : _GEN_5117; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5119 = 10'h2ff == io_inputs_1 ? 7'h0 : _GEN_5118; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5120 = 10'h300 == io_inputs_1 ? 7'h0 : _GEN_5119; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5121 = 10'h301 == io_inputs_1 ? 7'h0 : _GEN_5120; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5122 = 10'h302 == io_inputs_1 ? 7'h0 : _GEN_5121; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5123 = 10'h303 == io_inputs_1 ? 7'h0 : _GEN_5122; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5124 = 10'h304 == io_inputs_1 ? 7'h0 : _GEN_5123; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5125 = 10'h305 == io_inputs_1 ? 7'h0 : _GEN_5124; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5126 = 10'h306 == io_inputs_1 ? 7'h0 : _GEN_5125; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5127 = 10'h307 == io_inputs_1 ? 7'h0 : _GEN_5126; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5128 = 10'h308 == io_inputs_1 ? 7'h0 : _GEN_5127; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5129 = 10'h309 == io_inputs_1 ? 7'h0 : _GEN_5128; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5130 = 10'h30a == io_inputs_1 ? 7'h0 : _GEN_5129; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5131 = 10'h30b == io_inputs_1 ? 7'h0 : _GEN_5130; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5132 = 10'h30c == io_inputs_1 ? 7'h0 : _GEN_5131; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5133 = 10'h30d == io_inputs_1 ? 7'h0 : _GEN_5132; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5134 = 10'h30e == io_inputs_1 ? 7'h0 : _GEN_5133; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5135 = 10'h30f == io_inputs_1 ? 7'h0 : _GEN_5134; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5136 = 10'h310 == io_inputs_1 ? 7'h0 : _GEN_5135; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5137 = 10'h311 == io_inputs_1 ? 7'h0 : _GEN_5136; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5138 = 10'h312 == io_inputs_1 ? 7'h0 : _GEN_5137; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5139 = 10'h313 == io_inputs_1 ? 7'h0 : _GEN_5138; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5140 = 10'h314 == io_inputs_1 ? 7'h0 : _GEN_5139; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5141 = 10'h315 == io_inputs_1 ? 7'h0 : _GEN_5140; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5142 = 10'h316 == io_inputs_1 ? 7'h0 : _GEN_5141; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5143 = 10'h317 == io_inputs_1 ? 7'h0 : _GEN_5142; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5144 = 10'h318 == io_inputs_1 ? 7'h0 : _GEN_5143; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5145 = 10'h319 == io_inputs_1 ? 7'h0 : _GEN_5144; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5146 = 10'h31a == io_inputs_1 ? 7'h0 : _GEN_5145; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5147 = 10'h31b == io_inputs_1 ? 7'h0 : _GEN_5146; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5148 = 10'h31c == io_inputs_1 ? 7'h0 : _GEN_5147; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5149 = 10'h31d == io_inputs_1 ? 7'h0 : _GEN_5148; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5150 = 10'h31e == io_inputs_1 ? 7'h0 : _GEN_5149; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5151 = 10'h31f == io_inputs_1 ? 7'h0 : _GEN_5150; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5152 = 10'h320 == io_inputs_1 ? 7'h0 : _GEN_5151; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5153 = 10'h321 == io_inputs_1 ? 7'h0 : _GEN_5152; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5154 = 10'h322 == io_inputs_1 ? 7'h0 : _GEN_5153; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5155 = 10'h323 == io_inputs_1 ? 7'h0 : _GEN_5154; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5156 = 10'h324 == io_inputs_1 ? 7'h0 : _GEN_5155; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5157 = 10'h325 == io_inputs_1 ? 7'h0 : _GEN_5156; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5158 = 10'h326 == io_inputs_1 ? 7'h0 : _GEN_5157; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5159 = 10'h327 == io_inputs_1 ? 7'h0 : _GEN_5158; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5160 = 10'h328 == io_inputs_1 ? 7'h0 : _GEN_5159; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5161 = 10'h329 == io_inputs_1 ? 7'h0 : _GEN_5160; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5162 = 10'h32a == io_inputs_1 ? 7'h0 : _GEN_5161; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5163 = 10'h32b == io_inputs_1 ? 7'h0 : _GEN_5162; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5164 = 10'h32c == io_inputs_1 ? 7'h0 : _GEN_5163; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5165 = 10'h32d == io_inputs_1 ? 7'h0 : _GEN_5164; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5166 = 10'h32e == io_inputs_1 ? 7'h0 : _GEN_5165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5167 = 10'h32f == io_inputs_1 ? 7'h0 : _GEN_5166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5168 = 10'h330 == io_inputs_1 ? 7'h0 : _GEN_5167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5169 = 10'h331 == io_inputs_1 ? 7'h0 : _GEN_5168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5170 = 10'h332 == io_inputs_1 ? 7'h0 : _GEN_5169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5171 = 10'h333 == io_inputs_1 ? 7'h0 : _GEN_5170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5172 = 10'h334 == io_inputs_1 ? 7'h0 : _GEN_5171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5173 = 10'h335 == io_inputs_1 ? 7'h0 : _GEN_5172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5174 = 10'h336 == io_inputs_1 ? 7'h0 : _GEN_5173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5175 = 10'h337 == io_inputs_1 ? 7'h0 : _GEN_5174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5176 = 10'h338 == io_inputs_1 ? 7'h0 : _GEN_5175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5177 = 10'h339 == io_inputs_1 ? 7'h0 : _GEN_5176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5178 = 10'h33a == io_inputs_1 ? 7'h0 : _GEN_5177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5179 = 10'h33b == io_inputs_1 ? 7'h0 : _GEN_5178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5180 = 10'h33c == io_inputs_1 ? 7'h0 : _GEN_5179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5181 = 10'h33d == io_inputs_1 ? 7'h0 : _GEN_5180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5182 = 10'h33e == io_inputs_1 ? 7'h0 : _GEN_5181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5183 = 10'h33f == io_inputs_1 ? 7'h0 : _GEN_5182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5184 = 10'h340 == io_inputs_1 ? 7'h0 : _GEN_5183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5185 = 10'h341 == io_inputs_1 ? 7'h0 : _GEN_5184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5186 = 10'h342 == io_inputs_1 ? 7'h0 : _GEN_5185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5187 = 10'h343 == io_inputs_1 ? 7'h0 : _GEN_5186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5188 = 10'h344 == io_inputs_1 ? 7'h0 : _GEN_5187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5189 = 10'h345 == io_inputs_1 ? 7'h0 : _GEN_5188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5190 = 10'h346 == io_inputs_1 ? 7'h0 : _GEN_5189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5191 = 10'h347 == io_inputs_1 ? 7'h0 : _GEN_5190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5192 = 10'h348 == io_inputs_1 ? 7'h0 : _GEN_5191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5193 = 10'h349 == io_inputs_1 ? 7'h0 : _GEN_5192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5194 = 10'h34a == io_inputs_1 ? 7'h0 : _GEN_5193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5195 = 10'h34b == io_inputs_1 ? 7'h0 : _GEN_5194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5196 = 10'h34c == io_inputs_1 ? 7'h0 : _GEN_5195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5197 = 10'h34d == io_inputs_1 ? 7'h0 : _GEN_5196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5198 = 10'h34e == io_inputs_1 ? 7'h0 : _GEN_5197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5199 = 10'h34f == io_inputs_1 ? 7'h0 : _GEN_5198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5200 = 10'h350 == io_inputs_1 ? 7'h0 : _GEN_5199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5201 = 10'h351 == io_inputs_1 ? 7'h0 : _GEN_5200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5202 = 10'h352 == io_inputs_1 ? 7'h0 : _GEN_5201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5203 = 10'h353 == io_inputs_1 ? 7'h0 : _GEN_5202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5204 = 10'h354 == io_inputs_1 ? 7'h0 : _GEN_5203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5205 = 10'h355 == io_inputs_1 ? 7'h0 : _GEN_5204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5206 = 10'h356 == io_inputs_1 ? 7'h0 : _GEN_5205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5207 = 10'h357 == io_inputs_1 ? 7'h0 : _GEN_5206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5208 = 10'h358 == io_inputs_1 ? 7'h0 : _GEN_5207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5209 = 10'h359 == io_inputs_1 ? 7'h0 : _GEN_5208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5210 = 10'h35a == io_inputs_1 ? 7'h0 : _GEN_5209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5211 = 10'h35b == io_inputs_1 ? 7'h0 : _GEN_5210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5212 = 10'h35c == io_inputs_1 ? 7'h0 : _GEN_5211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5213 = 10'h35d == io_inputs_1 ? 7'h0 : _GEN_5212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5214 = 10'h35e == io_inputs_1 ? 7'h0 : _GEN_5213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5215 = 10'h35f == io_inputs_1 ? 7'h0 : _GEN_5214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5216 = 10'h360 == io_inputs_1 ? 7'h0 : _GEN_5215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5217 = 10'h361 == io_inputs_1 ? 7'h0 : _GEN_5216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5218 = 10'h362 == io_inputs_1 ? 7'h0 : _GEN_5217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5219 = 10'h363 == io_inputs_1 ? 7'h0 : _GEN_5218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5220 = 10'h364 == io_inputs_1 ? 7'h0 : _GEN_5219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5221 = 10'h365 == io_inputs_1 ? 7'h0 : _GEN_5220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5222 = 10'h366 == io_inputs_1 ? 7'h0 : _GEN_5221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5223 = 10'h367 == io_inputs_1 ? 7'h0 : _GEN_5222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5224 = 10'h368 == io_inputs_1 ? 7'h0 : _GEN_5223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5225 = 10'h369 == io_inputs_1 ? 7'h0 : _GEN_5224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5226 = 10'h36a == io_inputs_1 ? 7'h0 : _GEN_5225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5227 = 10'h36b == io_inputs_1 ? 7'h0 : _GEN_5226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5228 = 10'h36c == io_inputs_1 ? 7'h0 : _GEN_5227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5229 = 10'h36d == io_inputs_1 ? 7'h0 : _GEN_5228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5230 = 10'h36e == io_inputs_1 ? 7'h0 : _GEN_5229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5231 = 10'h36f == io_inputs_1 ? 7'h0 : _GEN_5230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5232 = 10'h370 == io_inputs_1 ? 7'h0 : _GEN_5231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5233 = 10'h371 == io_inputs_1 ? 7'h0 : _GEN_5232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5234 = 10'h372 == io_inputs_1 ? 7'h0 : _GEN_5233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5235 = 10'h373 == io_inputs_1 ? 7'h0 : _GEN_5234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5236 = 10'h374 == io_inputs_1 ? 7'h0 : _GEN_5235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5237 = 10'h375 == io_inputs_1 ? 7'h0 : _GEN_5236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5238 = 10'h376 == io_inputs_1 ? 7'h0 : _GEN_5237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5239 = 10'h377 == io_inputs_1 ? 7'h0 : _GEN_5238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5240 = 10'h378 == io_inputs_1 ? 7'h0 : _GEN_5239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5241 = 10'h379 == io_inputs_1 ? 7'h0 : _GEN_5240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5242 = 10'h37a == io_inputs_1 ? 7'h0 : _GEN_5241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5243 = 10'h37b == io_inputs_1 ? 7'h0 : _GEN_5242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5244 = 10'h37c == io_inputs_1 ? 7'h0 : _GEN_5243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5245 = 10'h37d == io_inputs_1 ? 7'h0 : _GEN_5244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5246 = 10'h37e == io_inputs_1 ? 7'h0 : _GEN_5245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5247 = 10'h37f == io_inputs_1 ? 7'h0 : _GEN_5246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5248 = 10'h380 == io_inputs_1 ? 7'h0 : _GEN_5247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5249 = 10'h381 == io_inputs_1 ? 7'h0 : _GEN_5248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5250 = 10'h382 == io_inputs_1 ? 7'h0 : _GEN_5249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5251 = 10'h383 == io_inputs_1 ? 7'h0 : _GEN_5250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5252 = 10'h384 == io_inputs_1 ? 7'h0 : _GEN_5251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5253 = 10'h385 == io_inputs_1 ? 7'h0 : _GEN_5252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5254 = 10'h386 == io_inputs_1 ? 7'h0 : _GEN_5253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5255 = 10'h387 == io_inputs_1 ? 7'h0 : _GEN_5254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5256 = 10'h388 == io_inputs_1 ? 7'h0 : _GEN_5255; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5257 = 10'h389 == io_inputs_1 ? 7'h0 : _GEN_5256; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5258 = 10'h38a == io_inputs_1 ? 7'h0 : _GEN_5257; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5259 = 10'h38b == io_inputs_1 ? 7'h0 : _GEN_5258; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5260 = 10'h38c == io_inputs_1 ? 7'h0 : _GEN_5259; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5261 = 10'h38d == io_inputs_1 ? 7'h0 : _GEN_5260; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5262 = 10'h38e == io_inputs_1 ? 7'h0 : _GEN_5261; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5263 = 10'h38f == io_inputs_1 ? 7'h0 : _GEN_5262; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5264 = 10'h390 == io_inputs_1 ? 7'h0 : _GEN_5263; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5265 = 10'h391 == io_inputs_1 ? 7'h0 : _GEN_5264; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5266 = 10'h392 == io_inputs_1 ? 7'h0 : _GEN_5265; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5267 = 10'h393 == io_inputs_1 ? 7'h0 : _GEN_5266; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5268 = 10'h394 == io_inputs_1 ? 7'h0 : _GEN_5267; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5269 = 10'h395 == io_inputs_1 ? 7'h0 : _GEN_5268; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5270 = 10'h396 == io_inputs_1 ? 7'h0 : _GEN_5269; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5271 = 10'h397 == io_inputs_1 ? 7'h0 : _GEN_5270; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5272 = 10'h398 == io_inputs_1 ? 7'h0 : _GEN_5271; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5273 = 10'h399 == io_inputs_1 ? 7'h0 : _GEN_5272; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5274 = 10'h39a == io_inputs_1 ? 7'h0 : _GEN_5273; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5275 = 10'h39b == io_inputs_1 ? 7'h0 : _GEN_5274; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5276 = 10'h39c == io_inputs_1 ? 7'h0 : _GEN_5275; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5277 = 10'h39d == io_inputs_1 ? 7'h0 : _GEN_5276; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5278 = 10'h39e == io_inputs_1 ? 7'h0 : _GEN_5277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5279 = 10'h39f == io_inputs_1 ? 7'h0 : _GEN_5278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5280 = 10'h3a0 == io_inputs_1 ? 7'h0 : _GEN_5279; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5281 = 10'h3a1 == io_inputs_1 ? 7'h0 : _GEN_5280; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5282 = 10'h3a2 == io_inputs_1 ? 7'h0 : _GEN_5281; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5283 = 10'h3a3 == io_inputs_1 ? 7'h0 : _GEN_5282; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5284 = 10'h3a4 == io_inputs_1 ? 7'h0 : _GEN_5283; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5285 = 10'h3a5 == io_inputs_1 ? 7'h0 : _GEN_5284; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5286 = 10'h3a6 == io_inputs_1 ? 7'h0 : _GEN_5285; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5287 = 10'h3a7 == io_inputs_1 ? 7'h0 : _GEN_5286; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5288 = 10'h3a8 == io_inputs_1 ? 7'h0 : _GEN_5287; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5289 = 10'h3a9 == io_inputs_1 ? 7'h0 : _GEN_5288; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5290 = 10'h3aa == io_inputs_1 ? 7'h0 : _GEN_5289; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5291 = 10'h3ab == io_inputs_1 ? 7'h0 : _GEN_5290; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5292 = 10'h3ac == io_inputs_1 ? 7'h0 : _GEN_5291; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5293 = 10'h3ad == io_inputs_1 ? 7'h0 : _GEN_5292; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5294 = 10'h3ae == io_inputs_1 ? 7'h0 : _GEN_5293; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5295 = 10'h3af == io_inputs_1 ? 7'h0 : _GEN_5294; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5296 = 10'h3b0 == io_inputs_1 ? 7'h0 : _GEN_5295; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5297 = 10'h3b1 == io_inputs_1 ? 7'h0 : _GEN_5296; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5298 = 10'h3b2 == io_inputs_1 ? 7'h0 : _GEN_5297; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5299 = 10'h3b3 == io_inputs_1 ? 7'h0 : _GEN_5298; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5300 = 10'h3b4 == io_inputs_1 ? 7'h0 : _GEN_5299; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5301 = 10'h3b5 == io_inputs_1 ? 7'h0 : _GEN_5300; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5302 = 10'h3b6 == io_inputs_1 ? 7'h0 : _GEN_5301; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5303 = 10'h3b7 == io_inputs_1 ? 7'h0 : _GEN_5302; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5304 = 10'h3b8 == io_inputs_1 ? 7'h0 : _GEN_5303; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5305 = 10'h3b9 == io_inputs_1 ? 7'h0 : _GEN_5304; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5306 = 10'h3ba == io_inputs_1 ? 7'h0 : _GEN_5305; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5307 = 10'h3bb == io_inputs_1 ? 7'h0 : _GEN_5306; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5308 = 10'h3bc == io_inputs_1 ? 7'h0 : _GEN_5307; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5309 = 10'h3bd == io_inputs_1 ? 7'h0 : _GEN_5308; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5310 = 10'h3be == io_inputs_1 ? 7'h0 : _GEN_5309; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5311 = 10'h3bf == io_inputs_1 ? 7'h0 : _GEN_5310; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5312 = 10'h3c0 == io_inputs_1 ? 7'h0 : _GEN_5311; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5313 = 10'h3c1 == io_inputs_1 ? 7'h0 : _GEN_5312; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5314 = 10'h3c2 == io_inputs_1 ? 7'h0 : _GEN_5313; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5315 = 10'h3c3 == io_inputs_1 ? 7'h0 : _GEN_5314; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5316 = 10'h3c4 == io_inputs_1 ? 7'h0 : _GEN_5315; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5317 = 10'h3c5 == io_inputs_1 ? 7'h0 : _GEN_5316; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5318 = 10'h3c6 == io_inputs_1 ? 7'h0 : _GEN_5317; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5319 = 10'h3c7 == io_inputs_1 ? 7'h0 : _GEN_5318; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5320 = 10'h3c8 == io_inputs_1 ? 7'h0 : _GEN_5319; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5321 = 10'h3c9 == io_inputs_1 ? 7'h0 : _GEN_5320; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5322 = 10'h3ca == io_inputs_1 ? 7'h0 : _GEN_5321; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5323 = 10'h3cb == io_inputs_1 ? 7'h0 : _GEN_5322; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5324 = 10'h3cc == io_inputs_1 ? 7'h0 : _GEN_5323; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5325 = 10'h3cd == io_inputs_1 ? 7'h0 : _GEN_5324; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5326 = 10'h3ce == io_inputs_1 ? 7'h0 : _GEN_5325; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5327 = 10'h3cf == io_inputs_1 ? 7'h0 : _GEN_5326; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5328 = 10'h3d0 == io_inputs_1 ? 7'h0 : _GEN_5327; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5329 = 10'h3d1 == io_inputs_1 ? 7'h0 : _GEN_5328; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5330 = 10'h3d2 == io_inputs_1 ? 7'h0 : _GEN_5329; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5331 = 10'h3d3 == io_inputs_1 ? 7'h0 : _GEN_5330; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5332 = 10'h3d4 == io_inputs_1 ? 7'h0 : _GEN_5331; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5333 = 10'h3d5 == io_inputs_1 ? 7'h0 : _GEN_5332; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5334 = 10'h3d6 == io_inputs_1 ? 7'h0 : _GEN_5333; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5335 = 10'h3d7 == io_inputs_1 ? 7'h0 : _GEN_5334; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5336 = 10'h3d8 == io_inputs_1 ? 7'h0 : _GEN_5335; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5337 = 10'h3d9 == io_inputs_1 ? 7'h0 : _GEN_5336; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5338 = 10'h3da == io_inputs_1 ? 7'h0 : _GEN_5337; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5339 = 10'h3db == io_inputs_1 ? 7'h0 : _GEN_5338; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5340 = 10'h3dc == io_inputs_1 ? 7'h0 : _GEN_5339; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5341 = 10'h3dd == io_inputs_1 ? 7'h0 : _GEN_5340; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5342 = 10'h3de == io_inputs_1 ? 7'h0 : _GEN_5341; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5343 = 10'h3df == io_inputs_1 ? 7'h0 : _GEN_5342; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5344 = 10'h3e0 == io_inputs_1 ? 7'h0 : _GEN_5343; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5345 = 10'h3e1 == io_inputs_1 ? 7'h0 : _GEN_5344; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5346 = 10'h3e2 == io_inputs_1 ? 7'h0 : _GEN_5345; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5347 = 10'h3e3 == io_inputs_1 ? 7'h0 : _GEN_5346; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5348 = 10'h3e4 == io_inputs_1 ? 7'h0 : _GEN_5347; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5349 = 10'h3e5 == io_inputs_1 ? 7'h0 : _GEN_5348; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5350 = 10'h3e6 == io_inputs_1 ? 7'h0 : _GEN_5349; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5351 = 10'h3e7 == io_inputs_1 ? 7'h0 : _GEN_5350; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5352 = 10'h3e8 == io_inputs_1 ? 7'h0 : _GEN_5351; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5353 = 10'h3e9 == io_inputs_1 ? 7'h0 : _GEN_5352; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5354 = 10'h3ea == io_inputs_1 ? 7'h0 : _GEN_5353; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5355 = 10'h3eb == io_inputs_1 ? 7'h0 : _GEN_5354; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5356 = 10'h3ec == io_inputs_1 ? 7'h0 : _GEN_5355; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5357 = 10'h3ed == io_inputs_1 ? 7'h0 : _GEN_5356; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5358 = 10'h3ee == io_inputs_1 ? 7'h0 : _GEN_5357; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5359 = 10'h3ef == io_inputs_1 ? 7'h0 : _GEN_5358; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5360 = 10'h3f0 == io_inputs_1 ? 7'h0 : _GEN_5359; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5361 = 10'h3f1 == io_inputs_1 ? 7'h0 : _GEN_5360; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5362 = 10'h3f2 == io_inputs_1 ? 7'h0 : _GEN_5361; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5363 = 10'h3f3 == io_inputs_1 ? 7'h0 : _GEN_5362; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5364 = 10'h3f4 == io_inputs_1 ? 7'h0 : _GEN_5363; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5365 = 10'h3f5 == io_inputs_1 ? 7'h0 : _GEN_5364; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5366 = 10'h3f6 == io_inputs_1 ? 7'h0 : _GEN_5365; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5367 = 10'h3f7 == io_inputs_1 ? 7'h0 : _GEN_5366; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5368 = 10'h3f8 == io_inputs_1 ? 7'h0 : _GEN_5367; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5369 = 10'h3f9 == io_inputs_1 ? 7'h0 : _GEN_5368; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5370 = 10'h3fa == io_inputs_1 ? 7'h0 : _GEN_5369; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5371 = 10'h3fb == io_inputs_1 ? 7'h0 : _GEN_5370; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5372 = 10'h3fc == io_inputs_1 ? 7'h0 : _GEN_5371; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5373 = 10'h3fd == io_inputs_1 ? 7'h0 : _GEN_5372; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5374 = 10'h3fe == io_inputs_1 ? 7'h0 : _GEN_5373; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5375 = 10'h3ff == io_inputs_1 ? 7'h0 : _GEN_5374; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5877 = 10'h1f5 == io_inputs_1 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5878 = 10'h1f6 == io_inputs_1 ? 7'h2 : _GEN_5877; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5879 = 10'h1f7 == io_inputs_1 ? 7'h3 : _GEN_5878; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5880 = 10'h1f8 == io_inputs_1 ? 7'h4 : _GEN_5879; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5881 = 10'h1f9 == io_inputs_1 ? 7'h5 : _GEN_5880; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5882 = 10'h1fa == io_inputs_1 ? 7'h6 : _GEN_5881; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5883 = 10'h1fb == io_inputs_1 ? 7'h7 : _GEN_5882; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5884 = 10'h1fc == io_inputs_1 ? 7'h8 : _GEN_5883; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5885 = 10'h1fd == io_inputs_1 ? 7'h9 : _GEN_5884; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5886 = 10'h1fe == io_inputs_1 ? 7'ha : _GEN_5885; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5887 = 10'h1ff == io_inputs_1 ? 7'hb : _GEN_5886; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5888 = 10'h200 == io_inputs_1 ? 7'hc : _GEN_5887; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5889 = 10'h201 == io_inputs_1 ? 7'hd : _GEN_5888; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5890 = 10'h202 == io_inputs_1 ? 7'he : _GEN_5889; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5891 = 10'h203 == io_inputs_1 ? 7'hf : _GEN_5890; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5892 = 10'h204 == io_inputs_1 ? 7'h10 : _GEN_5891; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5893 = 10'h205 == io_inputs_1 ? 7'h11 : _GEN_5892; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5894 = 10'h206 == io_inputs_1 ? 7'h12 : _GEN_5893; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5895 = 10'h207 == io_inputs_1 ? 7'h13 : _GEN_5894; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5896 = 10'h208 == io_inputs_1 ? 7'h14 : _GEN_5895; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5897 = 10'h209 == io_inputs_1 ? 7'h15 : _GEN_5896; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5898 = 10'h20a == io_inputs_1 ? 7'h16 : _GEN_5897; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5899 = 10'h20b == io_inputs_1 ? 7'h17 : _GEN_5898; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5900 = 10'h20c == io_inputs_1 ? 7'h18 : _GEN_5899; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5901 = 10'h20d == io_inputs_1 ? 7'h19 : _GEN_5900; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5902 = 10'h20e == io_inputs_1 ? 7'h1a : _GEN_5901; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5903 = 10'h20f == io_inputs_1 ? 7'h1b : _GEN_5902; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5904 = 10'h210 == io_inputs_1 ? 7'h1c : _GEN_5903; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5905 = 10'h211 == io_inputs_1 ? 7'h1d : _GEN_5904; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5906 = 10'h212 == io_inputs_1 ? 7'h1e : _GEN_5905; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5907 = 10'h213 == io_inputs_1 ? 7'h1f : _GEN_5906; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5908 = 10'h214 == io_inputs_1 ? 7'h20 : _GEN_5907; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5909 = 10'h215 == io_inputs_1 ? 7'h21 : _GEN_5908; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5910 = 10'h216 == io_inputs_1 ? 7'h22 : _GEN_5909; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5911 = 10'h217 == io_inputs_1 ? 7'h23 : _GEN_5910; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5912 = 10'h218 == io_inputs_1 ? 7'h24 : _GEN_5911; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5913 = 10'h219 == io_inputs_1 ? 7'h25 : _GEN_5912; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5914 = 10'h21a == io_inputs_1 ? 7'h26 : _GEN_5913; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5915 = 10'h21b == io_inputs_1 ? 7'h27 : _GEN_5914; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5916 = 10'h21c == io_inputs_1 ? 7'h28 : _GEN_5915; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5917 = 10'h21d == io_inputs_1 ? 7'h29 : _GEN_5916; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5918 = 10'h21e == io_inputs_1 ? 7'h2a : _GEN_5917; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5919 = 10'h21f == io_inputs_1 ? 7'h2b : _GEN_5918; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5920 = 10'h220 == io_inputs_1 ? 7'h2c : _GEN_5919; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5921 = 10'h221 == io_inputs_1 ? 7'h2d : _GEN_5920; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5922 = 10'h222 == io_inputs_1 ? 7'h2e : _GEN_5921; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5923 = 10'h223 == io_inputs_1 ? 7'h2f : _GEN_5922; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5924 = 10'h224 == io_inputs_1 ? 7'h30 : _GEN_5923; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5925 = 10'h225 == io_inputs_1 ? 7'h31 : _GEN_5924; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5926 = 10'h226 == io_inputs_1 ? 7'h32 : _GEN_5925; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5927 = 10'h227 == io_inputs_1 ? 7'h33 : _GEN_5926; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5928 = 10'h228 == io_inputs_1 ? 7'h34 : _GEN_5927; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5929 = 10'h229 == io_inputs_1 ? 7'h35 : _GEN_5928; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5930 = 10'h22a == io_inputs_1 ? 7'h36 : _GEN_5929; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5931 = 10'h22b == io_inputs_1 ? 7'h37 : _GEN_5930; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5932 = 10'h22c == io_inputs_1 ? 7'h38 : _GEN_5931; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5933 = 10'h22d == io_inputs_1 ? 7'h39 : _GEN_5932; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5934 = 10'h22e == io_inputs_1 ? 7'h3a : _GEN_5933; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5935 = 10'h22f == io_inputs_1 ? 7'h3b : _GEN_5934; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5936 = 10'h230 == io_inputs_1 ? 7'h3c : _GEN_5935; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5937 = 10'h231 == io_inputs_1 ? 7'h3d : _GEN_5936; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5938 = 10'h232 == io_inputs_1 ? 7'h3e : _GEN_5937; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5939 = 10'h233 == io_inputs_1 ? 7'h3f : _GEN_5938; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5940 = 10'h234 == io_inputs_1 ? 7'h40 : _GEN_5939; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5941 = 10'h235 == io_inputs_1 ? 7'h41 : _GEN_5940; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5942 = 10'h236 == io_inputs_1 ? 7'h42 : _GEN_5941; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5943 = 10'h237 == io_inputs_1 ? 7'h43 : _GEN_5942; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5944 = 10'h238 == io_inputs_1 ? 7'h44 : _GEN_5943; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5945 = 10'h239 == io_inputs_1 ? 7'h45 : _GEN_5944; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5946 = 10'h23a == io_inputs_1 ? 7'h46 : _GEN_5945; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5947 = 10'h23b == io_inputs_1 ? 7'h47 : _GEN_5946; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5948 = 10'h23c == io_inputs_1 ? 7'h48 : _GEN_5947; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5949 = 10'h23d == io_inputs_1 ? 7'h49 : _GEN_5948; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5950 = 10'h23e == io_inputs_1 ? 7'h4a : _GEN_5949; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5951 = 10'h23f == io_inputs_1 ? 7'h4b : _GEN_5950; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5952 = 10'h240 == io_inputs_1 ? 7'h4c : _GEN_5951; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5953 = 10'h241 == io_inputs_1 ? 7'h4d : _GEN_5952; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5954 = 10'h242 == io_inputs_1 ? 7'h4e : _GEN_5953; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5955 = 10'h243 == io_inputs_1 ? 7'h4f : _GEN_5954; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5956 = 10'h244 == io_inputs_1 ? 7'h50 : _GEN_5955; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5957 = 10'h245 == io_inputs_1 ? 7'h51 : _GEN_5956; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5958 = 10'h246 == io_inputs_1 ? 7'h52 : _GEN_5957; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5959 = 10'h247 == io_inputs_1 ? 7'h53 : _GEN_5958; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5960 = 10'h248 == io_inputs_1 ? 7'h54 : _GEN_5959; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5961 = 10'h249 == io_inputs_1 ? 7'h55 : _GEN_5960; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5962 = 10'h24a == io_inputs_1 ? 7'h56 : _GEN_5961; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5963 = 10'h24b == io_inputs_1 ? 7'h57 : _GEN_5962; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5964 = 10'h24c == io_inputs_1 ? 7'h58 : _GEN_5963; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5965 = 10'h24d == io_inputs_1 ? 7'h59 : _GEN_5964; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5966 = 10'h24e == io_inputs_1 ? 7'h5a : _GEN_5965; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5967 = 10'h24f == io_inputs_1 ? 7'h5b : _GEN_5966; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5968 = 10'h250 == io_inputs_1 ? 7'h5c : _GEN_5967; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5969 = 10'h251 == io_inputs_1 ? 7'h5d : _GEN_5968; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5970 = 10'h252 == io_inputs_1 ? 7'h5e : _GEN_5969; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5971 = 10'h253 == io_inputs_1 ? 7'h5f : _GEN_5970; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5972 = 10'h254 == io_inputs_1 ? 7'h60 : _GEN_5971; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5973 = 10'h255 == io_inputs_1 ? 7'h61 : _GEN_5972; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5974 = 10'h256 == io_inputs_1 ? 7'h62 : _GEN_5973; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5975 = 10'h257 == io_inputs_1 ? 7'h63 : _GEN_5974; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5976 = 10'h258 == io_inputs_1 ? 7'h64 : _GEN_5975; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5977 = 10'h259 == io_inputs_1 ? 7'h64 : _GEN_5976; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5978 = 10'h25a == io_inputs_1 ? 7'h64 : _GEN_5977; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5979 = 10'h25b == io_inputs_1 ? 7'h64 : _GEN_5978; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5980 = 10'h25c == io_inputs_1 ? 7'h64 : _GEN_5979; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5981 = 10'h25d == io_inputs_1 ? 7'h64 : _GEN_5980; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5982 = 10'h25e == io_inputs_1 ? 7'h64 : _GEN_5981; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5983 = 10'h25f == io_inputs_1 ? 7'h64 : _GEN_5982; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5984 = 10'h260 == io_inputs_1 ? 7'h64 : _GEN_5983; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5985 = 10'h261 == io_inputs_1 ? 7'h64 : _GEN_5984; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5986 = 10'h262 == io_inputs_1 ? 7'h64 : _GEN_5985; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5987 = 10'h263 == io_inputs_1 ? 7'h64 : _GEN_5986; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5988 = 10'h264 == io_inputs_1 ? 7'h64 : _GEN_5987; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5989 = 10'h265 == io_inputs_1 ? 7'h64 : _GEN_5988; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5990 = 10'h266 == io_inputs_1 ? 7'h64 : _GEN_5989; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5991 = 10'h267 == io_inputs_1 ? 7'h64 : _GEN_5990; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5992 = 10'h268 == io_inputs_1 ? 7'h64 : _GEN_5991; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5993 = 10'h269 == io_inputs_1 ? 7'h64 : _GEN_5992; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5994 = 10'h26a == io_inputs_1 ? 7'h64 : _GEN_5993; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5995 = 10'h26b == io_inputs_1 ? 7'h64 : _GEN_5994; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5996 = 10'h26c == io_inputs_1 ? 7'h64 : _GEN_5995; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5997 = 10'h26d == io_inputs_1 ? 7'h64 : _GEN_5996; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5998 = 10'h26e == io_inputs_1 ? 7'h64 : _GEN_5997; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_5999 = 10'h26f == io_inputs_1 ? 7'h64 : _GEN_5998; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6000 = 10'h270 == io_inputs_1 ? 7'h64 : _GEN_5999; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6001 = 10'h271 == io_inputs_1 ? 7'h64 : _GEN_6000; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6002 = 10'h272 == io_inputs_1 ? 7'h64 : _GEN_6001; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6003 = 10'h273 == io_inputs_1 ? 7'h64 : _GEN_6002; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6004 = 10'h274 == io_inputs_1 ? 7'h64 : _GEN_6003; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6005 = 10'h275 == io_inputs_1 ? 7'h64 : _GEN_6004; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6006 = 10'h276 == io_inputs_1 ? 7'h64 : _GEN_6005; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6007 = 10'h277 == io_inputs_1 ? 7'h64 : _GEN_6006; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6008 = 10'h278 == io_inputs_1 ? 7'h64 : _GEN_6007; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6009 = 10'h279 == io_inputs_1 ? 7'h64 : _GEN_6008; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6010 = 10'h27a == io_inputs_1 ? 7'h64 : _GEN_6009; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6011 = 10'h27b == io_inputs_1 ? 7'h64 : _GEN_6010; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6012 = 10'h27c == io_inputs_1 ? 7'h64 : _GEN_6011; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6013 = 10'h27d == io_inputs_1 ? 7'h64 : _GEN_6012; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6014 = 10'h27e == io_inputs_1 ? 7'h64 : _GEN_6013; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6015 = 10'h27f == io_inputs_1 ? 7'h64 : _GEN_6014; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6016 = 10'h280 == io_inputs_1 ? 7'h64 : _GEN_6015; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6017 = 10'h281 == io_inputs_1 ? 7'h64 : _GEN_6016; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6018 = 10'h282 == io_inputs_1 ? 7'h64 : _GEN_6017; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6019 = 10'h283 == io_inputs_1 ? 7'h64 : _GEN_6018; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6020 = 10'h284 == io_inputs_1 ? 7'h64 : _GEN_6019; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6021 = 10'h285 == io_inputs_1 ? 7'h64 : _GEN_6020; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6022 = 10'h286 == io_inputs_1 ? 7'h64 : _GEN_6021; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6023 = 10'h287 == io_inputs_1 ? 7'h64 : _GEN_6022; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6024 = 10'h288 == io_inputs_1 ? 7'h64 : _GEN_6023; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6025 = 10'h289 == io_inputs_1 ? 7'h64 : _GEN_6024; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6026 = 10'h28a == io_inputs_1 ? 7'h64 : _GEN_6025; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6027 = 10'h28b == io_inputs_1 ? 7'h64 : _GEN_6026; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6028 = 10'h28c == io_inputs_1 ? 7'h64 : _GEN_6027; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6029 = 10'h28d == io_inputs_1 ? 7'h64 : _GEN_6028; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6030 = 10'h28e == io_inputs_1 ? 7'h64 : _GEN_6029; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6031 = 10'h28f == io_inputs_1 ? 7'h64 : _GEN_6030; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6032 = 10'h290 == io_inputs_1 ? 7'h64 : _GEN_6031; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6033 = 10'h291 == io_inputs_1 ? 7'h64 : _GEN_6032; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6034 = 10'h292 == io_inputs_1 ? 7'h64 : _GEN_6033; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6035 = 10'h293 == io_inputs_1 ? 7'h64 : _GEN_6034; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6036 = 10'h294 == io_inputs_1 ? 7'h64 : _GEN_6035; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6037 = 10'h295 == io_inputs_1 ? 7'h64 : _GEN_6036; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6038 = 10'h296 == io_inputs_1 ? 7'h64 : _GEN_6037; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6039 = 10'h297 == io_inputs_1 ? 7'h64 : _GEN_6038; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6040 = 10'h298 == io_inputs_1 ? 7'h64 : _GEN_6039; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6041 = 10'h299 == io_inputs_1 ? 7'h64 : _GEN_6040; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6042 = 10'h29a == io_inputs_1 ? 7'h64 : _GEN_6041; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6043 = 10'h29b == io_inputs_1 ? 7'h64 : _GEN_6042; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6044 = 10'h29c == io_inputs_1 ? 7'h64 : _GEN_6043; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6045 = 10'h29d == io_inputs_1 ? 7'h64 : _GEN_6044; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6046 = 10'h29e == io_inputs_1 ? 7'h64 : _GEN_6045; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6047 = 10'h29f == io_inputs_1 ? 7'h64 : _GEN_6046; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6048 = 10'h2a0 == io_inputs_1 ? 7'h64 : _GEN_6047; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6049 = 10'h2a1 == io_inputs_1 ? 7'h64 : _GEN_6048; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6050 = 10'h2a2 == io_inputs_1 ? 7'h64 : _GEN_6049; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6051 = 10'h2a3 == io_inputs_1 ? 7'h64 : _GEN_6050; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6052 = 10'h2a4 == io_inputs_1 ? 7'h64 : _GEN_6051; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6053 = 10'h2a5 == io_inputs_1 ? 7'h64 : _GEN_6052; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6054 = 10'h2a6 == io_inputs_1 ? 7'h64 : _GEN_6053; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6055 = 10'h2a7 == io_inputs_1 ? 7'h64 : _GEN_6054; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6056 = 10'h2a8 == io_inputs_1 ? 7'h64 : _GEN_6055; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6057 = 10'h2a9 == io_inputs_1 ? 7'h64 : _GEN_6056; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6058 = 10'h2aa == io_inputs_1 ? 7'h64 : _GEN_6057; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6059 = 10'h2ab == io_inputs_1 ? 7'h64 : _GEN_6058; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6060 = 10'h2ac == io_inputs_1 ? 7'h64 : _GEN_6059; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6061 = 10'h2ad == io_inputs_1 ? 7'h64 : _GEN_6060; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6062 = 10'h2ae == io_inputs_1 ? 7'h64 : _GEN_6061; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6063 = 10'h2af == io_inputs_1 ? 7'h64 : _GEN_6062; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6064 = 10'h2b0 == io_inputs_1 ? 7'h64 : _GEN_6063; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6065 = 10'h2b1 == io_inputs_1 ? 7'h64 : _GEN_6064; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6066 = 10'h2b2 == io_inputs_1 ? 7'h64 : _GEN_6065; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6067 = 10'h2b3 == io_inputs_1 ? 7'h64 : _GEN_6066; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6068 = 10'h2b4 == io_inputs_1 ? 7'h64 : _GEN_6067; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6069 = 10'h2b5 == io_inputs_1 ? 7'h64 : _GEN_6068; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6070 = 10'h2b6 == io_inputs_1 ? 7'h64 : _GEN_6069; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6071 = 10'h2b7 == io_inputs_1 ? 7'h64 : _GEN_6070; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6072 = 10'h2b8 == io_inputs_1 ? 7'h64 : _GEN_6071; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6073 = 10'h2b9 == io_inputs_1 ? 7'h64 : _GEN_6072; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6074 = 10'h2ba == io_inputs_1 ? 7'h64 : _GEN_6073; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6075 = 10'h2bb == io_inputs_1 ? 7'h64 : _GEN_6074; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6076 = 10'h2bc == io_inputs_1 ? 7'h64 : _GEN_6075; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6077 = 10'h2bd == io_inputs_1 ? 7'h64 : _GEN_6076; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6078 = 10'h2be == io_inputs_1 ? 7'h64 : _GEN_6077; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6079 = 10'h2bf == io_inputs_1 ? 7'h64 : _GEN_6078; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6080 = 10'h2c0 == io_inputs_1 ? 7'h64 : _GEN_6079; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6081 = 10'h2c1 == io_inputs_1 ? 7'h64 : _GEN_6080; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6082 = 10'h2c2 == io_inputs_1 ? 7'h64 : _GEN_6081; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6083 = 10'h2c3 == io_inputs_1 ? 7'h64 : _GEN_6082; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6084 = 10'h2c4 == io_inputs_1 ? 7'h64 : _GEN_6083; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6085 = 10'h2c5 == io_inputs_1 ? 7'h64 : _GEN_6084; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6086 = 10'h2c6 == io_inputs_1 ? 7'h64 : _GEN_6085; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6087 = 10'h2c7 == io_inputs_1 ? 7'h64 : _GEN_6086; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6088 = 10'h2c8 == io_inputs_1 ? 7'h64 : _GEN_6087; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6089 = 10'h2c9 == io_inputs_1 ? 7'h64 : _GEN_6088; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6090 = 10'h2ca == io_inputs_1 ? 7'h64 : _GEN_6089; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6091 = 10'h2cb == io_inputs_1 ? 7'h64 : _GEN_6090; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6092 = 10'h2cc == io_inputs_1 ? 7'h64 : _GEN_6091; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6093 = 10'h2cd == io_inputs_1 ? 7'h64 : _GEN_6092; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6094 = 10'h2ce == io_inputs_1 ? 7'h64 : _GEN_6093; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6095 = 10'h2cf == io_inputs_1 ? 7'h64 : _GEN_6094; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6096 = 10'h2d0 == io_inputs_1 ? 7'h64 : _GEN_6095; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6097 = 10'h2d1 == io_inputs_1 ? 7'h64 : _GEN_6096; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6098 = 10'h2d2 == io_inputs_1 ? 7'h64 : _GEN_6097; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6099 = 10'h2d3 == io_inputs_1 ? 7'h64 : _GEN_6098; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6100 = 10'h2d4 == io_inputs_1 ? 7'h64 : _GEN_6099; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6101 = 10'h2d5 == io_inputs_1 ? 7'h64 : _GEN_6100; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6102 = 10'h2d6 == io_inputs_1 ? 7'h64 : _GEN_6101; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6103 = 10'h2d7 == io_inputs_1 ? 7'h64 : _GEN_6102; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6104 = 10'h2d8 == io_inputs_1 ? 7'h64 : _GEN_6103; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6105 = 10'h2d9 == io_inputs_1 ? 7'h64 : _GEN_6104; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6106 = 10'h2da == io_inputs_1 ? 7'h64 : _GEN_6105; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6107 = 10'h2db == io_inputs_1 ? 7'h64 : _GEN_6106; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6108 = 10'h2dc == io_inputs_1 ? 7'h64 : _GEN_6107; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6109 = 10'h2dd == io_inputs_1 ? 7'h64 : _GEN_6108; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6110 = 10'h2de == io_inputs_1 ? 7'h64 : _GEN_6109; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6111 = 10'h2df == io_inputs_1 ? 7'h64 : _GEN_6110; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6112 = 10'h2e0 == io_inputs_1 ? 7'h64 : _GEN_6111; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6113 = 10'h2e1 == io_inputs_1 ? 7'h64 : _GEN_6112; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6114 = 10'h2e2 == io_inputs_1 ? 7'h64 : _GEN_6113; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6115 = 10'h2e3 == io_inputs_1 ? 7'h64 : _GEN_6114; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6116 = 10'h2e4 == io_inputs_1 ? 7'h64 : _GEN_6115; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6117 = 10'h2e5 == io_inputs_1 ? 7'h64 : _GEN_6116; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6118 = 10'h2e6 == io_inputs_1 ? 7'h64 : _GEN_6117; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6119 = 10'h2e7 == io_inputs_1 ? 7'h64 : _GEN_6118; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6120 = 10'h2e8 == io_inputs_1 ? 7'h64 : _GEN_6119; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6121 = 10'h2e9 == io_inputs_1 ? 7'h64 : _GEN_6120; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6122 = 10'h2ea == io_inputs_1 ? 7'h64 : _GEN_6121; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6123 = 10'h2eb == io_inputs_1 ? 7'h64 : _GEN_6122; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6124 = 10'h2ec == io_inputs_1 ? 7'h64 : _GEN_6123; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6125 = 10'h2ed == io_inputs_1 ? 7'h64 : _GEN_6124; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6126 = 10'h2ee == io_inputs_1 ? 7'h64 : _GEN_6125; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6127 = 10'h2ef == io_inputs_1 ? 7'h64 : _GEN_6126; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6128 = 10'h2f0 == io_inputs_1 ? 7'h64 : _GEN_6127; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6129 = 10'h2f1 == io_inputs_1 ? 7'h64 : _GEN_6128; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6130 = 10'h2f2 == io_inputs_1 ? 7'h64 : _GEN_6129; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6131 = 10'h2f3 == io_inputs_1 ? 7'h64 : _GEN_6130; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6132 = 10'h2f4 == io_inputs_1 ? 7'h64 : _GEN_6131; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6133 = 10'h2f5 == io_inputs_1 ? 7'h64 : _GEN_6132; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6134 = 10'h2f6 == io_inputs_1 ? 7'h64 : _GEN_6133; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6135 = 10'h2f7 == io_inputs_1 ? 7'h64 : _GEN_6134; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6136 = 10'h2f8 == io_inputs_1 ? 7'h64 : _GEN_6135; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6137 = 10'h2f9 == io_inputs_1 ? 7'h64 : _GEN_6136; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6138 = 10'h2fa == io_inputs_1 ? 7'h64 : _GEN_6137; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6139 = 10'h2fb == io_inputs_1 ? 7'h64 : _GEN_6138; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6140 = 10'h2fc == io_inputs_1 ? 7'h64 : _GEN_6139; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6141 = 10'h2fd == io_inputs_1 ? 7'h64 : _GEN_6140; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6142 = 10'h2fe == io_inputs_1 ? 7'h64 : _GEN_6141; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6143 = 10'h2ff == io_inputs_1 ? 7'h64 : _GEN_6142; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6144 = 10'h300 == io_inputs_1 ? 7'h64 : _GEN_6143; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6145 = 10'h301 == io_inputs_1 ? 7'h64 : _GEN_6144; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6146 = 10'h302 == io_inputs_1 ? 7'h64 : _GEN_6145; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6147 = 10'h303 == io_inputs_1 ? 7'h64 : _GEN_6146; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6148 = 10'h304 == io_inputs_1 ? 7'h64 : _GEN_6147; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6149 = 10'h305 == io_inputs_1 ? 7'h64 : _GEN_6148; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6150 = 10'h306 == io_inputs_1 ? 7'h64 : _GEN_6149; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6151 = 10'h307 == io_inputs_1 ? 7'h64 : _GEN_6150; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6152 = 10'h308 == io_inputs_1 ? 7'h64 : _GEN_6151; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6153 = 10'h309 == io_inputs_1 ? 7'h64 : _GEN_6152; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6154 = 10'h30a == io_inputs_1 ? 7'h64 : _GEN_6153; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6155 = 10'h30b == io_inputs_1 ? 7'h64 : _GEN_6154; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6156 = 10'h30c == io_inputs_1 ? 7'h64 : _GEN_6155; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6157 = 10'h30d == io_inputs_1 ? 7'h64 : _GEN_6156; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6158 = 10'h30e == io_inputs_1 ? 7'h64 : _GEN_6157; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6159 = 10'h30f == io_inputs_1 ? 7'h64 : _GEN_6158; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6160 = 10'h310 == io_inputs_1 ? 7'h64 : _GEN_6159; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6161 = 10'h311 == io_inputs_1 ? 7'h64 : _GEN_6160; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6162 = 10'h312 == io_inputs_1 ? 7'h64 : _GEN_6161; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6163 = 10'h313 == io_inputs_1 ? 7'h64 : _GEN_6162; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6164 = 10'h314 == io_inputs_1 ? 7'h64 : _GEN_6163; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6165 = 10'h315 == io_inputs_1 ? 7'h64 : _GEN_6164; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6166 = 10'h316 == io_inputs_1 ? 7'h64 : _GEN_6165; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6167 = 10'h317 == io_inputs_1 ? 7'h64 : _GEN_6166; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6168 = 10'h318 == io_inputs_1 ? 7'h64 : _GEN_6167; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6169 = 10'h319 == io_inputs_1 ? 7'h64 : _GEN_6168; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6170 = 10'h31a == io_inputs_1 ? 7'h64 : _GEN_6169; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6171 = 10'h31b == io_inputs_1 ? 7'h64 : _GEN_6170; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6172 = 10'h31c == io_inputs_1 ? 7'h64 : _GEN_6171; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6173 = 10'h31d == io_inputs_1 ? 7'h64 : _GEN_6172; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6174 = 10'h31e == io_inputs_1 ? 7'h64 : _GEN_6173; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6175 = 10'h31f == io_inputs_1 ? 7'h64 : _GEN_6174; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6176 = 10'h320 == io_inputs_1 ? 7'h64 : _GEN_6175; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6177 = 10'h321 == io_inputs_1 ? 7'h64 : _GEN_6176; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6178 = 10'h322 == io_inputs_1 ? 7'h64 : _GEN_6177; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6179 = 10'h323 == io_inputs_1 ? 7'h64 : _GEN_6178; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6180 = 10'h324 == io_inputs_1 ? 7'h64 : _GEN_6179; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6181 = 10'h325 == io_inputs_1 ? 7'h64 : _GEN_6180; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6182 = 10'h326 == io_inputs_1 ? 7'h64 : _GEN_6181; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6183 = 10'h327 == io_inputs_1 ? 7'h64 : _GEN_6182; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6184 = 10'h328 == io_inputs_1 ? 7'h64 : _GEN_6183; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6185 = 10'h329 == io_inputs_1 ? 7'h64 : _GEN_6184; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6186 = 10'h32a == io_inputs_1 ? 7'h64 : _GEN_6185; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6187 = 10'h32b == io_inputs_1 ? 7'h64 : _GEN_6186; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6188 = 10'h32c == io_inputs_1 ? 7'h64 : _GEN_6187; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6189 = 10'h32d == io_inputs_1 ? 7'h64 : _GEN_6188; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6190 = 10'h32e == io_inputs_1 ? 7'h64 : _GEN_6189; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6191 = 10'h32f == io_inputs_1 ? 7'h64 : _GEN_6190; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6192 = 10'h330 == io_inputs_1 ? 7'h64 : _GEN_6191; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6193 = 10'h331 == io_inputs_1 ? 7'h64 : _GEN_6192; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6194 = 10'h332 == io_inputs_1 ? 7'h64 : _GEN_6193; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6195 = 10'h333 == io_inputs_1 ? 7'h64 : _GEN_6194; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6196 = 10'h334 == io_inputs_1 ? 7'h64 : _GEN_6195; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6197 = 10'h335 == io_inputs_1 ? 7'h64 : _GEN_6196; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6198 = 10'h336 == io_inputs_1 ? 7'h64 : _GEN_6197; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6199 = 10'h337 == io_inputs_1 ? 7'h64 : _GEN_6198; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6200 = 10'h338 == io_inputs_1 ? 7'h64 : _GEN_6199; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6201 = 10'h339 == io_inputs_1 ? 7'h64 : _GEN_6200; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6202 = 10'h33a == io_inputs_1 ? 7'h64 : _GEN_6201; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6203 = 10'h33b == io_inputs_1 ? 7'h64 : _GEN_6202; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6204 = 10'h33c == io_inputs_1 ? 7'h64 : _GEN_6203; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6205 = 10'h33d == io_inputs_1 ? 7'h64 : _GEN_6204; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6206 = 10'h33e == io_inputs_1 ? 7'h64 : _GEN_6205; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6207 = 10'h33f == io_inputs_1 ? 7'h64 : _GEN_6206; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6208 = 10'h340 == io_inputs_1 ? 7'h64 : _GEN_6207; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6209 = 10'h341 == io_inputs_1 ? 7'h64 : _GEN_6208; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6210 = 10'h342 == io_inputs_1 ? 7'h64 : _GEN_6209; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6211 = 10'h343 == io_inputs_1 ? 7'h64 : _GEN_6210; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6212 = 10'h344 == io_inputs_1 ? 7'h64 : _GEN_6211; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6213 = 10'h345 == io_inputs_1 ? 7'h64 : _GEN_6212; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6214 = 10'h346 == io_inputs_1 ? 7'h64 : _GEN_6213; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6215 = 10'h347 == io_inputs_1 ? 7'h64 : _GEN_6214; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6216 = 10'h348 == io_inputs_1 ? 7'h64 : _GEN_6215; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6217 = 10'h349 == io_inputs_1 ? 7'h64 : _GEN_6216; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6218 = 10'h34a == io_inputs_1 ? 7'h64 : _GEN_6217; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6219 = 10'h34b == io_inputs_1 ? 7'h64 : _GEN_6218; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6220 = 10'h34c == io_inputs_1 ? 7'h64 : _GEN_6219; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6221 = 10'h34d == io_inputs_1 ? 7'h64 : _GEN_6220; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6222 = 10'h34e == io_inputs_1 ? 7'h64 : _GEN_6221; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6223 = 10'h34f == io_inputs_1 ? 7'h64 : _GEN_6222; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6224 = 10'h350 == io_inputs_1 ? 7'h64 : _GEN_6223; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6225 = 10'h351 == io_inputs_1 ? 7'h64 : _GEN_6224; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6226 = 10'h352 == io_inputs_1 ? 7'h64 : _GEN_6225; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6227 = 10'h353 == io_inputs_1 ? 7'h64 : _GEN_6226; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6228 = 10'h354 == io_inputs_1 ? 7'h64 : _GEN_6227; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6229 = 10'h355 == io_inputs_1 ? 7'h64 : _GEN_6228; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6230 = 10'h356 == io_inputs_1 ? 7'h64 : _GEN_6229; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6231 = 10'h357 == io_inputs_1 ? 7'h64 : _GEN_6230; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6232 = 10'h358 == io_inputs_1 ? 7'h64 : _GEN_6231; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6233 = 10'h359 == io_inputs_1 ? 7'h64 : _GEN_6232; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6234 = 10'h35a == io_inputs_1 ? 7'h64 : _GEN_6233; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6235 = 10'h35b == io_inputs_1 ? 7'h64 : _GEN_6234; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6236 = 10'h35c == io_inputs_1 ? 7'h64 : _GEN_6235; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6237 = 10'h35d == io_inputs_1 ? 7'h64 : _GEN_6236; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6238 = 10'h35e == io_inputs_1 ? 7'h64 : _GEN_6237; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6239 = 10'h35f == io_inputs_1 ? 7'h64 : _GEN_6238; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6240 = 10'h360 == io_inputs_1 ? 7'h64 : _GEN_6239; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6241 = 10'h361 == io_inputs_1 ? 7'h64 : _GEN_6240; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6242 = 10'h362 == io_inputs_1 ? 7'h64 : _GEN_6241; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6243 = 10'h363 == io_inputs_1 ? 7'h64 : _GEN_6242; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6244 = 10'h364 == io_inputs_1 ? 7'h64 : _GEN_6243; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6245 = 10'h365 == io_inputs_1 ? 7'h64 : _GEN_6244; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6246 = 10'h366 == io_inputs_1 ? 7'h64 : _GEN_6245; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6247 = 10'h367 == io_inputs_1 ? 7'h64 : _GEN_6246; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6248 = 10'h368 == io_inputs_1 ? 7'h64 : _GEN_6247; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6249 = 10'h369 == io_inputs_1 ? 7'h64 : _GEN_6248; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6250 = 10'h36a == io_inputs_1 ? 7'h64 : _GEN_6249; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6251 = 10'h36b == io_inputs_1 ? 7'h64 : _GEN_6250; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6252 = 10'h36c == io_inputs_1 ? 7'h64 : _GEN_6251; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6253 = 10'h36d == io_inputs_1 ? 7'h64 : _GEN_6252; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6254 = 10'h36e == io_inputs_1 ? 7'h64 : _GEN_6253; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6255 = 10'h36f == io_inputs_1 ? 7'h64 : _GEN_6254; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6256 = 10'h370 == io_inputs_1 ? 7'h64 : _GEN_6255; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6257 = 10'h371 == io_inputs_1 ? 7'h64 : _GEN_6256; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6258 = 10'h372 == io_inputs_1 ? 7'h64 : _GEN_6257; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6259 = 10'h373 == io_inputs_1 ? 7'h64 : _GEN_6258; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6260 = 10'h374 == io_inputs_1 ? 7'h64 : _GEN_6259; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6261 = 10'h375 == io_inputs_1 ? 7'h64 : _GEN_6260; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6262 = 10'h376 == io_inputs_1 ? 7'h64 : _GEN_6261; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6263 = 10'h377 == io_inputs_1 ? 7'h64 : _GEN_6262; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6264 = 10'h378 == io_inputs_1 ? 7'h64 : _GEN_6263; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6265 = 10'h379 == io_inputs_1 ? 7'h64 : _GEN_6264; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6266 = 10'h37a == io_inputs_1 ? 7'h64 : _GEN_6265; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6267 = 10'h37b == io_inputs_1 ? 7'h64 : _GEN_6266; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6268 = 10'h37c == io_inputs_1 ? 7'h64 : _GEN_6267; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6269 = 10'h37d == io_inputs_1 ? 7'h64 : _GEN_6268; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6270 = 10'h37e == io_inputs_1 ? 7'h64 : _GEN_6269; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6271 = 10'h37f == io_inputs_1 ? 7'h64 : _GEN_6270; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6272 = 10'h380 == io_inputs_1 ? 7'h64 : _GEN_6271; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6273 = 10'h381 == io_inputs_1 ? 7'h64 : _GEN_6272; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6274 = 10'h382 == io_inputs_1 ? 7'h64 : _GEN_6273; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6275 = 10'h383 == io_inputs_1 ? 7'h64 : _GEN_6274; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6276 = 10'h384 == io_inputs_1 ? 7'h64 : _GEN_6275; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6277 = 10'h385 == io_inputs_1 ? 7'h64 : _GEN_6276; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6278 = 10'h386 == io_inputs_1 ? 7'h64 : _GEN_6277; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6279 = 10'h387 == io_inputs_1 ? 7'h64 : _GEN_6278; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6280 = 10'h388 == io_inputs_1 ? 7'h64 : _GEN_6279; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6281 = 10'h389 == io_inputs_1 ? 7'h64 : _GEN_6280; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6282 = 10'h38a == io_inputs_1 ? 7'h64 : _GEN_6281; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6283 = 10'h38b == io_inputs_1 ? 7'h64 : _GEN_6282; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6284 = 10'h38c == io_inputs_1 ? 7'h64 : _GEN_6283; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6285 = 10'h38d == io_inputs_1 ? 7'h64 : _GEN_6284; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6286 = 10'h38e == io_inputs_1 ? 7'h64 : _GEN_6285; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6287 = 10'h38f == io_inputs_1 ? 7'h64 : _GEN_6286; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6288 = 10'h390 == io_inputs_1 ? 7'h64 : _GEN_6287; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6289 = 10'h391 == io_inputs_1 ? 7'h64 : _GEN_6288; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6290 = 10'h392 == io_inputs_1 ? 7'h64 : _GEN_6289; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6291 = 10'h393 == io_inputs_1 ? 7'h64 : _GEN_6290; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6292 = 10'h394 == io_inputs_1 ? 7'h64 : _GEN_6291; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6293 = 10'h395 == io_inputs_1 ? 7'h64 : _GEN_6292; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6294 = 10'h396 == io_inputs_1 ? 7'h64 : _GEN_6293; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6295 = 10'h397 == io_inputs_1 ? 7'h64 : _GEN_6294; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6296 = 10'h398 == io_inputs_1 ? 7'h64 : _GEN_6295; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6297 = 10'h399 == io_inputs_1 ? 7'h64 : _GEN_6296; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6298 = 10'h39a == io_inputs_1 ? 7'h64 : _GEN_6297; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6299 = 10'h39b == io_inputs_1 ? 7'h64 : _GEN_6298; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6300 = 10'h39c == io_inputs_1 ? 7'h64 : _GEN_6299; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6301 = 10'h39d == io_inputs_1 ? 7'h64 : _GEN_6300; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6302 = 10'h39e == io_inputs_1 ? 7'h64 : _GEN_6301; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6303 = 10'h39f == io_inputs_1 ? 7'h64 : _GEN_6302; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6304 = 10'h3a0 == io_inputs_1 ? 7'h64 : _GEN_6303; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6305 = 10'h3a1 == io_inputs_1 ? 7'h64 : _GEN_6304; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6306 = 10'h3a2 == io_inputs_1 ? 7'h64 : _GEN_6305; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6307 = 10'h3a3 == io_inputs_1 ? 7'h64 : _GEN_6306; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6308 = 10'h3a4 == io_inputs_1 ? 7'h64 : _GEN_6307; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6309 = 10'h3a5 == io_inputs_1 ? 7'h64 : _GEN_6308; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6310 = 10'h3a6 == io_inputs_1 ? 7'h64 : _GEN_6309; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6311 = 10'h3a7 == io_inputs_1 ? 7'h64 : _GEN_6310; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6312 = 10'h3a8 == io_inputs_1 ? 7'h64 : _GEN_6311; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6313 = 10'h3a9 == io_inputs_1 ? 7'h64 : _GEN_6312; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6314 = 10'h3aa == io_inputs_1 ? 7'h64 : _GEN_6313; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6315 = 10'h3ab == io_inputs_1 ? 7'h64 : _GEN_6314; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6316 = 10'h3ac == io_inputs_1 ? 7'h64 : _GEN_6315; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6317 = 10'h3ad == io_inputs_1 ? 7'h64 : _GEN_6316; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6318 = 10'h3ae == io_inputs_1 ? 7'h64 : _GEN_6317; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6319 = 10'h3af == io_inputs_1 ? 7'h64 : _GEN_6318; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6320 = 10'h3b0 == io_inputs_1 ? 7'h64 : _GEN_6319; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6321 = 10'h3b1 == io_inputs_1 ? 7'h64 : _GEN_6320; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6322 = 10'h3b2 == io_inputs_1 ? 7'h64 : _GEN_6321; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6323 = 10'h3b3 == io_inputs_1 ? 7'h64 : _GEN_6322; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6324 = 10'h3b4 == io_inputs_1 ? 7'h64 : _GEN_6323; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6325 = 10'h3b5 == io_inputs_1 ? 7'h64 : _GEN_6324; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6326 = 10'h3b6 == io_inputs_1 ? 7'h64 : _GEN_6325; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6327 = 10'h3b7 == io_inputs_1 ? 7'h64 : _GEN_6326; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6328 = 10'h3b8 == io_inputs_1 ? 7'h64 : _GEN_6327; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6329 = 10'h3b9 == io_inputs_1 ? 7'h64 : _GEN_6328; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6330 = 10'h3ba == io_inputs_1 ? 7'h64 : _GEN_6329; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6331 = 10'h3bb == io_inputs_1 ? 7'h64 : _GEN_6330; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6332 = 10'h3bc == io_inputs_1 ? 7'h64 : _GEN_6331; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6333 = 10'h3bd == io_inputs_1 ? 7'h64 : _GEN_6332; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6334 = 10'h3be == io_inputs_1 ? 7'h64 : _GEN_6333; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6335 = 10'h3bf == io_inputs_1 ? 7'h64 : _GEN_6334; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6336 = 10'h3c0 == io_inputs_1 ? 7'h64 : _GEN_6335; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6337 = 10'h3c1 == io_inputs_1 ? 7'h64 : _GEN_6336; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6338 = 10'h3c2 == io_inputs_1 ? 7'h64 : _GEN_6337; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6339 = 10'h3c3 == io_inputs_1 ? 7'h64 : _GEN_6338; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6340 = 10'h3c4 == io_inputs_1 ? 7'h64 : _GEN_6339; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6341 = 10'h3c5 == io_inputs_1 ? 7'h64 : _GEN_6340; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6342 = 10'h3c6 == io_inputs_1 ? 7'h64 : _GEN_6341; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6343 = 10'h3c7 == io_inputs_1 ? 7'h64 : _GEN_6342; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6344 = 10'h3c8 == io_inputs_1 ? 7'h64 : _GEN_6343; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6345 = 10'h3c9 == io_inputs_1 ? 7'h64 : _GEN_6344; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6346 = 10'h3ca == io_inputs_1 ? 7'h64 : _GEN_6345; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6347 = 10'h3cb == io_inputs_1 ? 7'h64 : _GEN_6346; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6348 = 10'h3cc == io_inputs_1 ? 7'h64 : _GEN_6347; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6349 = 10'h3cd == io_inputs_1 ? 7'h64 : _GEN_6348; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6350 = 10'h3ce == io_inputs_1 ? 7'h64 : _GEN_6349; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6351 = 10'h3cf == io_inputs_1 ? 7'h64 : _GEN_6350; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6352 = 10'h3d0 == io_inputs_1 ? 7'h64 : _GEN_6351; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6353 = 10'h3d1 == io_inputs_1 ? 7'h64 : _GEN_6352; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6354 = 10'h3d2 == io_inputs_1 ? 7'h64 : _GEN_6353; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6355 = 10'h3d3 == io_inputs_1 ? 7'h64 : _GEN_6354; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6356 = 10'h3d4 == io_inputs_1 ? 7'h64 : _GEN_6355; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6357 = 10'h3d5 == io_inputs_1 ? 7'h64 : _GEN_6356; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6358 = 10'h3d6 == io_inputs_1 ? 7'h64 : _GEN_6357; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6359 = 10'h3d7 == io_inputs_1 ? 7'h64 : _GEN_6358; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6360 = 10'h3d8 == io_inputs_1 ? 7'h64 : _GEN_6359; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6361 = 10'h3d9 == io_inputs_1 ? 7'h64 : _GEN_6360; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6362 = 10'h3da == io_inputs_1 ? 7'h64 : _GEN_6361; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6363 = 10'h3db == io_inputs_1 ? 7'h64 : _GEN_6362; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6364 = 10'h3dc == io_inputs_1 ? 7'h64 : _GEN_6363; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6365 = 10'h3dd == io_inputs_1 ? 7'h64 : _GEN_6364; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6366 = 10'h3de == io_inputs_1 ? 7'h64 : _GEN_6365; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6367 = 10'h3df == io_inputs_1 ? 7'h64 : _GEN_6366; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6368 = 10'h3e0 == io_inputs_1 ? 7'h64 : _GEN_6367; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6369 = 10'h3e1 == io_inputs_1 ? 7'h64 : _GEN_6368; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6370 = 10'h3e2 == io_inputs_1 ? 7'h64 : _GEN_6369; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6371 = 10'h3e3 == io_inputs_1 ? 7'h64 : _GEN_6370; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6372 = 10'h3e4 == io_inputs_1 ? 7'h64 : _GEN_6371; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6373 = 10'h3e5 == io_inputs_1 ? 7'h64 : _GEN_6372; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6374 = 10'h3e6 == io_inputs_1 ? 7'h64 : _GEN_6373; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6375 = 10'h3e7 == io_inputs_1 ? 7'h64 : _GEN_6374; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6376 = 10'h3e8 == io_inputs_1 ? 7'h64 : _GEN_6375; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6377 = 10'h3e9 == io_inputs_1 ? 7'h64 : _GEN_6376; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6378 = 10'h3ea == io_inputs_1 ? 7'h64 : _GEN_6377; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6379 = 10'h3eb == io_inputs_1 ? 7'h64 : _GEN_6378; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6380 = 10'h3ec == io_inputs_1 ? 7'h64 : _GEN_6379; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6381 = 10'h3ed == io_inputs_1 ? 7'h64 : _GEN_6380; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6382 = 10'h3ee == io_inputs_1 ? 7'h64 : _GEN_6381; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6383 = 10'h3ef == io_inputs_1 ? 7'h64 : _GEN_6382; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6384 = 10'h3f0 == io_inputs_1 ? 7'h64 : _GEN_6383; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6385 = 10'h3f1 == io_inputs_1 ? 7'h64 : _GEN_6384; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6386 = 10'h3f2 == io_inputs_1 ? 7'h64 : _GEN_6385; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6387 = 10'h3f3 == io_inputs_1 ? 7'h64 : _GEN_6386; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6388 = 10'h3f4 == io_inputs_1 ? 7'h64 : _GEN_6387; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6389 = 10'h3f5 == io_inputs_1 ? 7'h64 : _GEN_6388; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6390 = 10'h3f6 == io_inputs_1 ? 7'h64 : _GEN_6389; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6391 = 10'h3f7 == io_inputs_1 ? 7'h64 : _GEN_6390; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6392 = 10'h3f8 == io_inputs_1 ? 7'h64 : _GEN_6391; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6393 = 10'h3f9 == io_inputs_1 ? 7'h64 : _GEN_6392; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6394 = 10'h3fa == io_inputs_1 ? 7'h64 : _GEN_6393; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6395 = 10'h3fb == io_inputs_1 ? 7'h64 : _GEN_6394; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6396 = 10'h3fc == io_inputs_1 ? 7'h64 : _GEN_6395; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6397 = 10'h3fd == io_inputs_1 ? 7'h64 : _GEN_6396; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6398 = 10'h3fe == io_inputs_1 ? 7'h64 : _GEN_6397; // @[regular_fuzzification.scala 177:{36,36}]
  wire [6:0] _GEN_6399 = 10'h3ff == io_inputs_1 ? 7'h64 : _GEN_6398; // @[regular_fuzzification.scala 177:{36,36}]
  wire  regMinVec_0_maxMinOutput = regMinVec_0_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_1_maxMinOutput = regMinVec_1_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_2_maxMinOutput = regMinVec_2_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_3_maxMinOutput = regMinVec_3_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_4_maxMinOutput = regMinVec_4_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_5_maxMinOutput = regMinVec_5_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_6_maxMinOutput = regMinVec_6_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_7_maxMinOutput = regMinVec_7_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_8_maxMinOutput = regMinVec_8_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_9_maxMinOutput = regMinVec_9_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_10_maxMinOutput = regMinVec_10_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_11_maxMinOutput = regMinVec_11_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_12_maxMinOutput = regMinVec_12_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_13_maxMinOutput = regMinVec_13_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_14_maxMinOutput = regMinVec_14_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_15_maxMinOutput = regMinVec_15_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_16_maxMinOutput = regMinVec_16_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_17_maxMinOutput = regMinVec_17_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_18_maxMinOutput = regMinVec_18_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_19_maxMinOutput = regMinVec_19_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_20_maxMinOutput = regMinVec_20_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_21_maxMinOutput = regMinVec_21_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_22_maxMinOutput = regMinVec_22_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_23_maxMinOutput = regMinVec_23_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_24_maxMinOutput = regMinVec_24_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire [6:0] _GEN_6425 = io_start ? _GEN_255 : {{4'd0}, regLutResultsVec_0}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6426 = io_start ? _GEN_511 : {{4'd0}, regLutResultsVec_1}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6427 = io_start ? _GEN_767 : {{4'd0}, regLutResultsVec_2}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6428 = io_start ? _GEN_1023 : {{4'd0}, regLutResultsVec_3}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6429 = io_start ? _GEN_1279 : {{4'd0}, regLutResultsVec_4}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6430 = io_start ? _GEN_2303 : {{4'd0}, regLutResultsVec_5}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6431 = io_start ? _GEN_3327 : {{4'd0}, regLutResultsVec_6}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6432 = io_start ? _GEN_4351 : {{4'd0}, regLutResultsVec_7}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6433 = io_start ? _GEN_5375 : {{4'd0}, regLutResultsVec_8}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [6:0] _GEN_6434 = io_start ? _GEN_6399 : {{4'd0}, regLutResultsVec_9}; // @[regular_fuzzification.scala 125:29 164:29 177:36]
  wire [2:0] regMaxVec_0_result = regMaxVec_0_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_1_result = regMaxVec_1_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_2_result = regMaxVec_2_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_3_result = regMaxVec_3_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_4_result = regMaxVec_4_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] outResult_result = outResult_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  Comparator regMinVec_0_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_0_comparatorModule_io_in1),
    .io_in2(regMinVec_0_comparatorModule_io_in2),
    .io_maxMin(regMinVec_0_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_1_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_1_comparatorModule_io_in1),
    .io_in2(regMinVec_1_comparatorModule_io_in2),
    .io_maxMin(regMinVec_1_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_2_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_2_comparatorModule_io_in1),
    .io_in2(regMinVec_2_comparatorModule_io_in2),
    .io_maxMin(regMinVec_2_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_3_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_3_comparatorModule_io_in1),
    .io_in2(regMinVec_3_comparatorModule_io_in2),
    .io_maxMin(regMinVec_3_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_4_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_4_comparatorModule_io_in1),
    .io_in2(regMinVec_4_comparatorModule_io_in2),
    .io_maxMin(regMinVec_4_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_5_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_5_comparatorModule_io_in1),
    .io_in2(regMinVec_5_comparatorModule_io_in2),
    .io_maxMin(regMinVec_5_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_6_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_6_comparatorModule_io_in1),
    .io_in2(regMinVec_6_comparatorModule_io_in2),
    .io_maxMin(regMinVec_6_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_7_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_7_comparatorModule_io_in1),
    .io_in2(regMinVec_7_comparatorModule_io_in2),
    .io_maxMin(regMinVec_7_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_8_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_8_comparatorModule_io_in1),
    .io_in2(regMinVec_8_comparatorModule_io_in2),
    .io_maxMin(regMinVec_8_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_9_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_9_comparatorModule_io_in1),
    .io_in2(regMinVec_9_comparatorModule_io_in2),
    .io_maxMin(regMinVec_9_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_10_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_10_comparatorModule_io_in1),
    .io_in2(regMinVec_10_comparatorModule_io_in2),
    .io_maxMin(regMinVec_10_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_11_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_11_comparatorModule_io_in1),
    .io_in2(regMinVec_11_comparatorModule_io_in2),
    .io_maxMin(regMinVec_11_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_12_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_12_comparatorModule_io_in1),
    .io_in2(regMinVec_12_comparatorModule_io_in2),
    .io_maxMin(regMinVec_12_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_13_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_13_comparatorModule_io_in1),
    .io_in2(regMinVec_13_comparatorModule_io_in2),
    .io_maxMin(regMinVec_13_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_14_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_14_comparatorModule_io_in1),
    .io_in2(regMinVec_14_comparatorModule_io_in2),
    .io_maxMin(regMinVec_14_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_15_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_15_comparatorModule_io_in1),
    .io_in2(regMinVec_15_comparatorModule_io_in2),
    .io_maxMin(regMinVec_15_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_16_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_16_comparatorModule_io_in1),
    .io_in2(regMinVec_16_comparatorModule_io_in2),
    .io_maxMin(regMinVec_16_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_17_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_17_comparatorModule_io_in1),
    .io_in2(regMinVec_17_comparatorModule_io_in2),
    .io_maxMin(regMinVec_17_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_18_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_18_comparatorModule_io_in1),
    .io_in2(regMinVec_18_comparatorModule_io_in2),
    .io_maxMin(regMinVec_18_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_19_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_19_comparatorModule_io_in1),
    .io_in2(regMinVec_19_comparatorModule_io_in2),
    .io_maxMin(regMinVec_19_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_20_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_20_comparatorModule_io_in1),
    .io_in2(regMinVec_20_comparatorModule_io_in2),
    .io_maxMin(regMinVec_20_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_21_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_21_comparatorModule_io_in1),
    .io_in2(regMinVec_21_comparatorModule_io_in2),
    .io_maxMin(regMinVec_21_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_22_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_22_comparatorModule_io_in1),
    .io_in2(regMinVec_22_comparatorModule_io_in2),
    .io_maxMin(regMinVec_22_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_23_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_23_comparatorModule_io_in1),
    .io_in2(regMinVec_23_comparatorModule_io_in2),
    .io_maxMin(regMinVec_23_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_24_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_24_comparatorModule_io_in1),
    .io_in2(regMinVec_24_comparatorModule_io_in2),
    .io_maxMin(regMinVec_24_comparatorModule_io_maxMin)
  );
  MultipleComparator regMaxVec_0_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_0_comparatorModule_clock),
    .io_start(regMaxVec_0_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_0_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_0_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_0_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_0_comparatorModule_io_inputs_3),
    .io_result(regMaxVec_0_comparatorModule_io_result)
  );
  MultipleComparator_1 regMaxVec_1_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_1_comparatorModule_clock),
    .io_start(regMaxVec_1_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_1_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_1_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_1_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_1_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_1_comparatorModule_io_inputs_4),
    .io_inputs_5(regMaxVec_1_comparatorModule_io_inputs_5),
    .io_result(regMaxVec_1_comparatorModule_io_result)
  );
  MultipleComparator regMaxVec_2_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_2_comparatorModule_clock),
    .io_start(regMaxVec_2_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_2_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_2_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_2_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_2_comparatorModule_io_inputs_3),
    .io_result(regMaxVec_2_comparatorModule_io_result)
  );
  MultipleComparator_1 regMaxVec_3_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_3_comparatorModule_clock),
    .io_start(regMaxVec_3_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_3_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_3_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_3_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_3_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_3_comparatorModule_io_inputs_4),
    .io_inputs_5(regMaxVec_3_comparatorModule_io_inputs_5),
    .io_result(regMaxVec_3_comparatorModule_io_result)
  );
  MultipleComparator_4 regMaxVec_4_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_4_comparatorModule_clock),
    .io_start(regMaxVec_4_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_4_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_4_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_4_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_4_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_4_comparatorModule_io_inputs_4),
    .io_result(regMaxVec_4_comparatorModule_io_result)
  );
  MultipleComparator_5 outResult_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(outResult_comparatorModule_clock),
    .io_start(outResult_comparatorModule_io_start),
    .io_inputs_0(outResult_comparatorModule_io_inputs_0),
    .io_inputs_1(outResult_comparatorModule_io_inputs_1),
    .io_inputs_2(outResult_comparatorModule_io_inputs_2),
    .io_inputs_3(outResult_comparatorModule_io_inputs_3),
    .io_inputs_4(outResult_comparatorModule_io_inputs_4),
    .io_result(outResult_comparatorModule_io_result)
  );
  assign io_outResultValid = 1'h0; // @[regular_fuzzification.scala 164:29 399:20]
  assign io_outResult = io_start ? outResult_result : 3'h0; // @[regular_fuzzification.scala 164:29 373:15 398:15]
  assign regMinVec_0_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_0_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_1_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_1_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_2_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_2_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_3_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_3_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_4_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_4_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_5_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_5_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_6_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_6_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_7_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_7_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_8_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_8_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_9_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_9_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_10_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_10_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_11_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_11_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_12_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_12_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_13_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_13_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_14_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_14_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_15_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_15_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_16_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_16_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_17_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_17_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_18_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_18_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_19_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_19_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_20_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_20_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_21_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_21_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_22_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_22_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_23_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_23_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_24_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_24_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMaxVec_0_comparatorModule_clock = clock;
  assign regMaxVec_0_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_0_comparatorModule_io_inputs_0 = regMinVec_0; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_0_comparatorModule_io_inputs_1 = regMinVec_1; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_0_comparatorModule_io_inputs_2 = regMinVec_2; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_0_comparatorModule_io_inputs_3 = regMinVec_5; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_1_comparatorModule_clock = clock;
  assign regMaxVec_1_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_1_comparatorModule_io_inputs_0 = regMinVec_3; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_1_comparatorModule_io_inputs_1 = regMinVec_4; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_1_comparatorModule_io_inputs_2 = regMinVec_6; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_1_comparatorModule_io_inputs_3 = regMinVec_7; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_1_comparatorModule_io_inputs_4 = regMinVec_8; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_1_comparatorModule_io_inputs_5 = regMinVec_10; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_2_comparatorModule_clock = clock;
  assign regMaxVec_2_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_2_comparatorModule_io_inputs_0 = regMinVec_9; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_2_comparatorModule_io_inputs_1 = regMinVec_11; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_2_comparatorModule_io_inputs_2 = regMinVec_12; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_2_comparatorModule_io_inputs_3 = regMinVec_15; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_3_comparatorModule_clock = clock;
  assign regMaxVec_3_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_3_comparatorModule_io_inputs_0 = regMinVec_13; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_3_comparatorModule_io_inputs_1 = regMinVec_14; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_3_comparatorModule_io_inputs_2 = regMinVec_16; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_3_comparatorModule_io_inputs_3 = regMinVec_17; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_3_comparatorModule_io_inputs_4 = regMinVec_20; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_3_comparatorModule_io_inputs_5 = regMinVec_21; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_4_comparatorModule_clock = clock;
  assign regMaxVec_4_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_4_comparatorModule_io_inputs_0 = regMinVec_18; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_4_comparatorModule_io_inputs_1 = regMinVec_19; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_4_comparatorModule_io_inputs_2 = regMinVec_22; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_4_comparatorModule_io_inputs_3 = regMinVec_23; // @[regular_fuzzification.scala 301:15 304:30]
  assign regMaxVec_4_comparatorModule_io_inputs_4 = regMinVec_24; // @[regular_fuzzification.scala 301:15 304:30]
  assign outResult_comparatorModule_clock = clock;
  assign outResult_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign outResult_comparatorModule_io_inputs_0 = regMaxVec_0; // @[regular_fuzzification.scala 356:11 363:40]
  assign outResult_comparatorModule_io_inputs_1 = regMaxVec_1; // @[regular_fuzzification.scala 356:11 363:40]
  assign outResult_comparatorModule_io_inputs_2 = regMaxVec_2; // @[regular_fuzzification.scala 356:11 363:40]
  assign outResult_comparatorModule_io_inputs_3 = regMaxVec_3; // @[regular_fuzzification.scala 356:11 363:40]
  assign outResult_comparatorModule_io_inputs_4 = regMaxVec_4; // @[regular_fuzzification.scala 356:11 363:40]
  always @(posedge clock) begin
    regLutResultsVec_0 <= _GEN_6425[2:0];
    regLutResultsVec_1 <= _GEN_6426[2:0];
    regLutResultsVec_2 <= _GEN_6427[2:0];
    regLutResultsVec_3 <= _GEN_6428[2:0];
    regLutResultsVec_4 <= _GEN_6429[2:0];
    regLutResultsVec_5 <= _GEN_6430[2:0];
    regLutResultsVec_6 <= _GEN_6431[2:0];
    regLutResultsVec_7 <= _GEN_6432[2:0];
    regLutResultsVec_8 <= _GEN_6433[2:0];
    regLutResultsVec_9 <= _GEN_6434[2:0];
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_0_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_0 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_0 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_1_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_1 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_1 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_2_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_2 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_2 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_3_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_3 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_3 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_4_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_4 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_4 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_5_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_5 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_5 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_6_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_6 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_6 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_7_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_7 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_7 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_8_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_8 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_8 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_9_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_9 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_9 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_10_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_10 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_10 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_11_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_11 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_11 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_12_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_12 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_12 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_13_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_13 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_13 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_14_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_14 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_14 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_15_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_15 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_15 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_16_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_16 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_16 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_17_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_17 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_17 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_18_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_18 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_18 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_19_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_19 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_19 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_20_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_20 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_20 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_21_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_21 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_21 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_22_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_22 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_22 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_23_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_23 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_23 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      if (~regMinVec_24_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_24 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_24 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      regMaxVec_0 <= regMaxVec_0_result; // @[regular_fuzzification.scala 307:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      regMaxVec_1 <= regMaxVec_1_result; // @[regular_fuzzification.scala 307:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      regMaxVec_2 <= regMaxVec_2_result; // @[regular_fuzzification.scala 307:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      regMaxVec_3 <= regMaxVec_3_result; // @[regular_fuzzification.scala 307:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 164:29]
      regMaxVec_4 <= regMaxVec_4_result; // @[regular_fuzzification.scala 307:39]
    end
  end
endmodule
