module LutMembershipFunctionOnline_1(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [9:0] i; // @[lut_mem_online.scala 215:18]
  reg  buffer_0; // @[lut_mem_online.scala 219:19]
  reg  buffer_1; // @[lut_mem_online.scala 219:19]
  reg  buffer_2; // @[lut_mem_online.scala 219:19]
  reg  buffer_3; // @[lut_mem_online.scala 219:19]
  reg  buffer_4; // @[lut_mem_online.scala 219:19]
  reg  buffer_5; // @[lut_mem_online.scala 219:19]
  reg  buffer_6; // @[lut_mem_online.scala 219:19]
  reg [4:0] counter; // @[lut_mem_online.scala 221:24]
  reg  outResult; // @[lut_mem_online.scala 224:26]
  wire  _T_2 = counter < 5'ha; // @[lut_mem_online.scala 241:22]
  wire  _GEN_0 = io_inputBit ? 1'h0 : buffer_0; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_1 = i == 10'h0 ? _GEN_0 : buffer_0; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_2 = io_inputBit ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_3 = i == 10'h1 ? _GEN_2 : _GEN_1; // @[lut_mem_online.scala 247:34]
  wire  _GEN_4 = io_inputBit ? 1'h0 : _GEN_3; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_5 = i == 10'h3 ? _GEN_4 : _GEN_3; // @[lut_mem_online.scala 247:34]
  wire  _T_10 = ~io_inputBit; // @[lut_mem_online.scala 249:32]
  wire  _GEN_6 = ~io_inputBit | _GEN_5; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_7 = i == 10'h7 ? _GEN_6 : _GEN_5; // @[lut_mem_online.scala 247:34]
  wire  _GEN_8 = io_inputBit ? 1'h0 : _GEN_7; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_9 = i == 10'h10 ? _GEN_8 : _GEN_7; // @[lut_mem_online.scala 247:34]
  wire  _GEN_10 = ~io_inputBit | _GEN_9; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_11 = i == 10'h21 ? _GEN_10 : _GEN_9; // @[lut_mem_online.scala 247:34]
  wire  _GEN_12 = io_inputBit ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_13 = i == 10'h44 ? _GEN_12 : _GEN_11; // @[lut_mem_online.scala 247:34]
  wire  _GEN_14 = ~io_inputBit | _GEN_13; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_15 = i == 10'h89 ? _GEN_14 : _GEN_13; // @[lut_mem_online.scala 247:34]
  wire  _GEN_16 = ~io_inputBit | _GEN_15; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_17 = i == 10'h114 ? _GEN_16 : _GEN_15; // @[lut_mem_online.scala 247:34]
  wire  _GEN_18 = ~io_inputBit | _GEN_17; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_19 = i == 10'h22a ? _GEN_18 : _GEN_17; // @[lut_mem_online.scala 247:34]
  wire  _GEN_20 = io_inputBit ? 1'h0 : _GEN_19; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_21 = i == 10'h22a ? _GEN_20 : _GEN_19; // @[lut_mem_online.scala 247:34]
  wire  _GEN_22 = io_inputBit ? 1'h0 : buffer_1; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_23 = i == 10'h0 ? _GEN_22 : buffer_1; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_24 = io_inputBit ? 1'h0 : _GEN_23; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_25 = i == 10'h1 ? _GEN_24 : _GEN_23; // @[lut_mem_online.scala 247:34]
  wire  _GEN_26 = io_inputBit ? 1'h0 : _GEN_25; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_27 = i == 10'h3 ? _GEN_26 : _GEN_25; // @[lut_mem_online.scala 247:34]
  wire  _GEN_28 = ~io_inputBit | _GEN_27; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_29 = i == 10'hf ? _GEN_28 : _GEN_27; // @[lut_mem_online.scala 247:34]
  wire  _GEN_30 = ~io_inputBit | _GEN_29; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_31 = i == 10'h20 ? _GEN_30 : _GEN_29; // @[lut_mem_online.scala 247:34]
  wire  _GEN_32 = ~io_inputBit ? 1'h0 : _GEN_31; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_33 = i == 10'h21 ? _GEN_32 : _GEN_31; // @[lut_mem_online.scala 247:34]
  wire  _GEN_34 = ~io_inputBit | _GEN_33; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_35 = i == 10'h22 ? _GEN_34 : _GEN_33; // @[lut_mem_online.scala 247:34]
  wire  _GEN_36 = io_inputBit ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_37 = i == 10'h42 ? _GEN_36 : _GEN_35; // @[lut_mem_online.scala 247:34]
  wire  _GEN_38 = io_inputBit | _GEN_37; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_39 = i == 10'h44 ? _GEN_38 : _GEN_37; // @[lut_mem_online.scala 247:34]
  wire  _GEN_40 = io_inputBit ? 1'h0 : _GEN_39; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_41 = i == 10'h46 ? _GEN_40 : _GEN_39; // @[lut_mem_online.scala 247:34]
  wire  _GEN_42 = ~io_inputBit | _GEN_41; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_43 = i == 10'h85 ? _GEN_42 : _GEN_41; // @[lut_mem_online.scala 247:34]
  wire  _GEN_44 = ~io_inputBit ? 1'h0 : _GEN_43; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_45 = i == 10'h89 ? _GEN_44 : _GEN_43; // @[lut_mem_online.scala 247:34]
  wire  _GEN_46 = ~io_inputBit | _GEN_45; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_47 = i == 10'h8d ? _GEN_46 : _GEN_45; // @[lut_mem_online.scala 247:34]
  wire  _GEN_48 = ~io_inputBit | _GEN_47; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_49 = i == 10'h10c ? _GEN_48 : _GEN_47; // @[lut_mem_online.scala 247:34]
  wire  _GEN_50 = ~io_inputBit ? 1'h0 : _GEN_49; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_51 = i == 10'h114 ? _GEN_50 : _GEN_49; // @[lut_mem_online.scala 247:34]
  wire  _GEN_52 = ~io_inputBit | _GEN_51; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_53 = i == 10'h11c ? _GEN_52 : _GEN_51; // @[lut_mem_online.scala 247:34]
  wire  _GEN_54 = ~io_inputBit | _GEN_53; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_55 = i == 10'h21a ? _GEN_54 : _GEN_53; // @[lut_mem_online.scala 247:34]
  wire  _GEN_56 = io_inputBit ? 1'h0 : _GEN_55; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_57 = i == 10'h21a ? _GEN_56 : _GEN_55; // @[lut_mem_online.scala 247:34]
  wire  _GEN_58 = ~io_inputBit ? 1'h0 : _GEN_57; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_59 = i == 10'h22a ? _GEN_58 : _GEN_57; // @[lut_mem_online.scala 247:34]
  wire  _GEN_60 = io_inputBit | _GEN_59; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_61 = i == 10'h22a ? _GEN_60 : _GEN_59; // @[lut_mem_online.scala 247:34]
  wire  _GEN_62 = ~io_inputBit | _GEN_61; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_63 = i == 10'h23a ? _GEN_62 : _GEN_61; // @[lut_mem_online.scala 247:34]
  wire  _GEN_64 = io_inputBit ? 1'h0 : _GEN_63; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_65 = i == 10'h23a ? _GEN_64 : _GEN_63; // @[lut_mem_online.scala 247:34]
  wire  _GEN_66 = io_inputBit ? 1'h0 : buffer_2; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_67 = i == 10'h0 ? _GEN_66 : buffer_2; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_68 = io_inputBit ? 1'h0 : _GEN_67; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_69 = i == 10'h1 ? _GEN_68 : _GEN_67; // @[lut_mem_online.scala 247:34]
  wire  _GEN_70 = io_inputBit ? 1'h0 : _GEN_69; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_71 = i == 10'h8 ? _GEN_70 : _GEN_69; // @[lut_mem_online.scala 247:34]
  wire  _GEN_72 = ~io_inputBit ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_73 = i == 10'hf ? _GEN_72 : _GEN_71; // @[lut_mem_online.scala 247:34]
  wire  _GEN_74 = io_inputBit ? 1'h0 : _GEN_73; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_75 = i == 10'h11 ? _GEN_74 : _GEN_73; // @[lut_mem_online.scala 247:34]
  wire  _GEN_76 = ~io_inputBit ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_77 = i == 10'h20 ? _GEN_76 : _GEN_75; // @[lut_mem_online.scala 247:34]
  wire  _GEN_78 = io_inputBit ? 1'h0 : _GEN_77; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_79 = i == 10'h23 ? _GEN_78 : _GEN_77; // @[lut_mem_online.scala 247:34]
  wire  _GEN_80 = io_inputBit | _GEN_79; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_81 = i == 10'h42 ? _GEN_80 : _GEN_79; // @[lut_mem_online.scala 247:34]
  wire  _GEN_82 = io_inputBit ? 1'h0 : _GEN_81; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_83 = i == 10'h43 ? _GEN_82 : _GEN_81; // @[lut_mem_online.scala 247:34]
  wire  _GEN_84 = io_inputBit | _GEN_83; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_85 = i == 10'h44 ? _GEN_84 : _GEN_83; // @[lut_mem_online.scala 247:34]
  wire  _GEN_86 = io_inputBit ? 1'h0 : _GEN_85; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_87 = i == 10'h45 ? _GEN_86 : _GEN_85; // @[lut_mem_online.scala 247:34]
  wire  _GEN_88 = io_inputBit | _GEN_87; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_89 = i == 10'h46 ? _GEN_88 : _GEN_87; // @[lut_mem_online.scala 247:34]
  wire  _GEN_90 = io_inputBit ? 1'h0 : _GEN_89; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_91 = i == 10'h47 ? _GEN_90 : _GEN_89; // @[lut_mem_online.scala 247:34]
  wire  _GEN_92 = ~io_inputBit ? 1'h0 : _GEN_91; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_93 = i == 10'h85 ? _GEN_92 : _GEN_91; // @[lut_mem_online.scala 247:34]
  wire  _GEN_94 = ~io_inputBit | _GEN_93; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_95 = i == 10'h87 ? _GEN_94 : _GEN_93; // @[lut_mem_online.scala 247:34]
  wire  _GEN_96 = ~io_inputBit ? 1'h0 : _GEN_95; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_97 = i == 10'h89 ? _GEN_96 : _GEN_95; // @[lut_mem_online.scala 247:34]
  wire  _GEN_98 = ~io_inputBit | _GEN_97; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_99 = i == 10'h8b ? _GEN_98 : _GEN_97; // @[lut_mem_online.scala 247:34]
  wire  _GEN_100 = ~io_inputBit ? 1'h0 : _GEN_99; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_101 = i == 10'h8d ? _GEN_100 : _GEN_99; // @[lut_mem_online.scala 247:34]
  wire  _GEN_102 = ~io_inputBit | _GEN_101; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_103 = i == 10'h8f ? _GEN_102 : _GEN_101; // @[lut_mem_online.scala 247:34]
  wire  _GEN_104 = ~io_inputBit ? 1'h0 : _GEN_103; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_105 = i == 10'h10c ? _GEN_104 : _GEN_103; // @[lut_mem_online.scala 247:34]
  wire  _GEN_106 = ~io_inputBit | _GEN_105; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_107 = i == 10'h110 ? _GEN_106 : _GEN_105; // @[lut_mem_online.scala 247:34]
  wire  _GEN_108 = ~io_inputBit ? 1'h0 : _GEN_107; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_109 = i == 10'h114 ? _GEN_108 : _GEN_107; // @[lut_mem_online.scala 247:34]
  wire  _GEN_110 = ~io_inputBit | _GEN_109; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_111 = i == 10'h118 ? _GEN_110 : _GEN_109; // @[lut_mem_online.scala 247:34]
  wire  _GEN_112 = ~io_inputBit ? 1'h0 : _GEN_111; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_113 = i == 10'h11c ? _GEN_112 : _GEN_111; // @[lut_mem_online.scala 247:34]
  wire  _GEN_114 = ~io_inputBit | _GEN_113; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_115 = i == 10'h120 ? _GEN_114 : _GEN_113; // @[lut_mem_online.scala 247:34]
  wire  _GEN_116 = ~io_inputBit ? 1'h0 : _GEN_115; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_117 = i == 10'h21a ? _GEN_116 : _GEN_115; // @[lut_mem_online.scala 247:34]
  wire  _GEN_118 = io_inputBit | _GEN_117; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_119 = i == 10'h21a ? _GEN_118 : _GEN_117; // @[lut_mem_online.scala 247:34]
  wire  _GEN_120 = ~io_inputBit | _GEN_119; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_121 = i == 10'h222 ? _GEN_120 : _GEN_119; // @[lut_mem_online.scala 247:34]
  wire  _GEN_122 = io_inputBit ? 1'h0 : _GEN_121; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_123 = i == 10'h222 ? _GEN_122 : _GEN_121; // @[lut_mem_online.scala 247:34]
  wire  _GEN_124 = ~io_inputBit ? 1'h0 : _GEN_123; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_125 = i == 10'h22a ? _GEN_124 : _GEN_123; // @[lut_mem_online.scala 247:34]
  wire  _GEN_126 = io_inputBit | _GEN_125; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_127 = i == 10'h22a ? _GEN_126 : _GEN_125; // @[lut_mem_online.scala 247:34]
  wire  _GEN_128 = ~io_inputBit | _GEN_127; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_129 = i == 10'h232 ? _GEN_128 : _GEN_127; // @[lut_mem_online.scala 247:34]
  wire  _GEN_130 = io_inputBit ? 1'h0 : _GEN_129; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_131 = i == 10'h232 ? _GEN_130 : _GEN_129; // @[lut_mem_online.scala 247:34]
  wire  _GEN_132 = ~io_inputBit ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_133 = i == 10'h23a ? _GEN_132 : _GEN_131; // @[lut_mem_online.scala 247:34]
  wire  _GEN_134 = io_inputBit | _GEN_133; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_135 = i == 10'h23a ? _GEN_134 : _GEN_133; // @[lut_mem_online.scala 247:34]
  wire  _GEN_136 = ~io_inputBit | _GEN_135; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_137 = i == 10'h242 ? _GEN_136 : _GEN_135; // @[lut_mem_online.scala 247:34]
  wire  _GEN_138 = io_inputBit ? 1'h0 : _GEN_137; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_139 = i == 10'h242 ? _GEN_138 : _GEN_137; // @[lut_mem_online.scala 247:34]
  wire  _GEN_140 = io_inputBit ? 1'h0 : buffer_3; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_141 = i == 10'h0 ? _GEN_140 : buffer_3; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_142 = io_inputBit ? 1'h0 : _GEN_141; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_143 = i == 10'h1 ? _GEN_142 : _GEN_141; // @[lut_mem_online.scala 247:34]
  wire  _GEN_144 = io_inputBit ? 1'h0 : _GEN_143; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_145 = i == 10'h8 ? _GEN_144 : _GEN_143; // @[lut_mem_online.scala 247:34]
  wire  _GEN_146 = ~io_inputBit ? 1'h0 : _GEN_145; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_147 = i == 10'hf ? _GEN_146 : _GEN_145; // @[lut_mem_online.scala 247:34]
  wire  _GEN_148 = io_inputBit ? 1'h0 : _GEN_147; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_149 = i == 10'h11 ? _GEN_148 : _GEN_147; // @[lut_mem_online.scala 247:34]
  wire  _GEN_150 = ~io_inputBit ? 1'h0 : _GEN_149; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_151 = i == 10'h20 ? _GEN_150 : _GEN_149; // @[lut_mem_online.scala 247:34]
  wire  _GEN_152 = io_inputBit ? 1'h0 : _GEN_151; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_153 = i == 10'h23 ? _GEN_152 : _GEN_151; // @[lut_mem_online.scala 247:34]
  wire  _GEN_154 = ~io_inputBit ? 1'h0 : _GEN_153; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_155 = i == 10'h85 ? _GEN_154 : _GEN_153; // @[lut_mem_online.scala 247:34]
  wire  _GEN_156 = ~io_inputBit | _GEN_155; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_157 = i == 10'h86 ? _GEN_156 : _GEN_155; // @[lut_mem_online.scala 247:34]
  wire  _GEN_158 = ~io_inputBit ? 1'h0 : _GEN_157; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_159 = i == 10'h87 ? _GEN_158 : _GEN_157; // @[lut_mem_online.scala 247:34]
  wire  _GEN_160 = ~io_inputBit | _GEN_159; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_161 = i == 10'h88 ? _GEN_160 : _GEN_159; // @[lut_mem_online.scala 247:34]
  wire  _GEN_162 = ~io_inputBit ? 1'h0 : _GEN_161; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_163 = i == 10'h89 ? _GEN_162 : _GEN_161; // @[lut_mem_online.scala 247:34]
  wire  _GEN_164 = ~io_inputBit | _GEN_163; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_165 = i == 10'h8a ? _GEN_164 : _GEN_163; // @[lut_mem_online.scala 247:34]
  wire  _GEN_166 = ~io_inputBit ? 1'h0 : _GEN_165; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_167 = i == 10'h8b ? _GEN_166 : _GEN_165; // @[lut_mem_online.scala 247:34]
  wire  _GEN_168 = ~io_inputBit | _GEN_167; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_169 = i == 10'h8c ? _GEN_168 : _GEN_167; // @[lut_mem_online.scala 247:34]
  wire  _GEN_170 = ~io_inputBit ? 1'h0 : _GEN_169; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_171 = i == 10'h8d ? _GEN_170 : _GEN_169; // @[lut_mem_online.scala 247:34]
  wire  _GEN_172 = ~io_inputBit | _GEN_171; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_173 = i == 10'h8e ? _GEN_172 : _GEN_171; // @[lut_mem_online.scala 247:34]
  wire  _GEN_174 = ~io_inputBit ? 1'h0 : _GEN_173; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_175 = i == 10'h8f ? _GEN_174 : _GEN_173; // @[lut_mem_online.scala 247:34]
  wire  _GEN_176 = ~io_inputBit | _GEN_175; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_177 = i == 10'h90 ? _GEN_176 : _GEN_175; // @[lut_mem_online.scala 247:34]
  wire  _GEN_178 = ~io_inputBit ? 1'h0 : _GEN_177; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_179 = i == 10'h10c ? _GEN_178 : _GEN_177; // @[lut_mem_online.scala 247:34]
  wire  _GEN_180 = ~io_inputBit | _GEN_179; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_181 = i == 10'h10e ? _GEN_180 : _GEN_179; // @[lut_mem_online.scala 247:34]
  wire  _GEN_182 = ~io_inputBit ? 1'h0 : _GEN_181; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_183 = i == 10'h110 ? _GEN_182 : _GEN_181; // @[lut_mem_online.scala 247:34]
  wire  _GEN_184 = ~io_inputBit | _GEN_183; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_185 = i == 10'h112 ? _GEN_184 : _GEN_183; // @[lut_mem_online.scala 247:34]
  wire  _GEN_186 = ~io_inputBit ? 1'h0 : _GEN_185; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_187 = i == 10'h114 ? _GEN_186 : _GEN_185; // @[lut_mem_online.scala 247:34]
  wire  _GEN_188 = ~io_inputBit | _GEN_187; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_189 = i == 10'h116 ? _GEN_188 : _GEN_187; // @[lut_mem_online.scala 247:34]
  wire  _GEN_190 = ~io_inputBit ? 1'h0 : _GEN_189; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_191 = i == 10'h118 ? _GEN_190 : _GEN_189; // @[lut_mem_online.scala 247:34]
  wire  _GEN_192 = ~io_inputBit | _GEN_191; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_193 = i == 10'h11a ? _GEN_192 : _GEN_191; // @[lut_mem_online.scala 247:34]
  wire  _GEN_194 = ~io_inputBit ? 1'h0 : _GEN_193; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_195 = i == 10'h11c ? _GEN_194 : _GEN_193; // @[lut_mem_online.scala 247:34]
  wire  _GEN_196 = ~io_inputBit | _GEN_195; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_197 = i == 10'h11e ? _GEN_196 : _GEN_195; // @[lut_mem_online.scala 247:34]
  wire  _GEN_198 = ~io_inputBit ? 1'h0 : _GEN_197; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_199 = i == 10'h120 ? _GEN_198 : _GEN_197; // @[lut_mem_online.scala 247:34]
  wire  _GEN_200 = ~io_inputBit | _GEN_199; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_201 = i == 10'h122 ? _GEN_200 : _GEN_199; // @[lut_mem_online.scala 247:34]
  wire  _GEN_202 = ~io_inputBit ? 1'h0 : _GEN_201; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_203 = i == 10'h21a ? _GEN_202 : _GEN_201; // @[lut_mem_online.scala 247:34]
  wire  _GEN_204 = io_inputBit | _GEN_203; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_205 = i == 10'h21a ? _GEN_204 : _GEN_203; // @[lut_mem_online.scala 247:34]
  wire  _GEN_206 = ~io_inputBit | _GEN_205; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_207 = i == 10'h21e ? _GEN_206 : _GEN_205; // @[lut_mem_online.scala 247:34]
  wire  _GEN_208 = io_inputBit ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_209 = i == 10'h21e ? _GEN_208 : _GEN_207; // @[lut_mem_online.scala 247:34]
  wire  _GEN_210 = ~io_inputBit ? 1'h0 : _GEN_209; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_211 = i == 10'h222 ? _GEN_210 : _GEN_209; // @[lut_mem_online.scala 247:34]
  wire  _GEN_212 = io_inputBit | _GEN_211; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_213 = i == 10'h222 ? _GEN_212 : _GEN_211; // @[lut_mem_online.scala 247:34]
  wire  _GEN_214 = ~io_inputBit | _GEN_213; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_215 = i == 10'h226 ? _GEN_214 : _GEN_213; // @[lut_mem_online.scala 247:34]
  wire  _GEN_216 = io_inputBit ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_217 = i == 10'h226 ? _GEN_216 : _GEN_215; // @[lut_mem_online.scala 247:34]
  wire  _GEN_218 = ~io_inputBit ? 1'h0 : _GEN_217; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_219 = i == 10'h22a ? _GEN_218 : _GEN_217; // @[lut_mem_online.scala 247:34]
  wire  _GEN_220 = io_inputBit | _GEN_219; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_221 = i == 10'h22a ? _GEN_220 : _GEN_219; // @[lut_mem_online.scala 247:34]
  wire  _GEN_222 = ~io_inputBit | _GEN_221; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_223 = i == 10'h22e ? _GEN_222 : _GEN_221; // @[lut_mem_online.scala 247:34]
  wire  _GEN_224 = io_inputBit ? 1'h0 : _GEN_223; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_225 = i == 10'h22e ? _GEN_224 : _GEN_223; // @[lut_mem_online.scala 247:34]
  wire  _GEN_226 = ~io_inputBit ? 1'h0 : _GEN_225; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_227 = i == 10'h232 ? _GEN_226 : _GEN_225; // @[lut_mem_online.scala 247:34]
  wire  _GEN_228 = io_inputBit | _GEN_227; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_229 = i == 10'h232 ? _GEN_228 : _GEN_227; // @[lut_mem_online.scala 247:34]
  wire  _GEN_230 = ~io_inputBit | _GEN_229; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_231 = i == 10'h236 ? _GEN_230 : _GEN_229; // @[lut_mem_online.scala 247:34]
  wire  _GEN_232 = io_inputBit ? 1'h0 : _GEN_231; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_233 = i == 10'h236 ? _GEN_232 : _GEN_231; // @[lut_mem_online.scala 247:34]
  wire  _GEN_234 = ~io_inputBit ? 1'h0 : _GEN_233; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_235 = i == 10'h23a ? _GEN_234 : _GEN_233; // @[lut_mem_online.scala 247:34]
  wire  _GEN_236 = io_inputBit | _GEN_235; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_237 = i == 10'h23a ? _GEN_236 : _GEN_235; // @[lut_mem_online.scala 247:34]
  wire  _GEN_238 = ~io_inputBit | _GEN_237; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_239 = i == 10'h23e ? _GEN_238 : _GEN_237; // @[lut_mem_online.scala 247:34]
  wire  _GEN_240 = io_inputBit ? 1'h0 : _GEN_239; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_241 = i == 10'h23e ? _GEN_240 : _GEN_239; // @[lut_mem_online.scala 247:34]
  wire  _GEN_242 = ~io_inputBit ? 1'h0 : _GEN_241; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_243 = i == 10'h242 ? _GEN_242 : _GEN_241; // @[lut_mem_online.scala 247:34]
  wire  _GEN_244 = io_inputBit | _GEN_243; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_245 = i == 10'h242 ? _GEN_244 : _GEN_243; // @[lut_mem_online.scala 247:34]
  wire  _GEN_246 = ~io_inputBit | _GEN_245; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_247 = i == 10'h246 ? _GEN_246 : _GEN_245; // @[lut_mem_online.scala 247:34]
  wire  _GEN_248 = io_inputBit ? 1'h0 : _GEN_247; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_249 = i == 10'h246 ? _GEN_248 : _GEN_247; // @[lut_mem_online.scala 247:34]
  wire  _GEN_250 = io_inputBit ? 1'h0 : buffer_4; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_251 = i == 10'h0 ? _GEN_250 : buffer_4; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_252 = io_inputBit ? 1'h0 : _GEN_251; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_253 = i == 10'h1 ? _GEN_252 : _GEN_251; // @[lut_mem_online.scala 247:34]
  wire  _GEN_254 = io_inputBit ? 1'h0 : _GEN_253; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_255 = i == 10'h8 ? _GEN_254 : _GEN_253; // @[lut_mem_online.scala 247:34]
  wire  _GEN_256 = ~io_inputBit | _GEN_255; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_257 = i == 10'hf ? _GEN_256 : _GEN_255; // @[lut_mem_online.scala 247:34]
  wire  _GEN_258 = io_inputBit ? 1'h0 : _GEN_257; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_259 = i == 10'h11 ? _GEN_258 : _GEN_257; // @[lut_mem_online.scala 247:34]
  wire  _GEN_260 = ~io_inputBit | _GEN_259; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_261 = i == 10'h20 ? _GEN_260 : _GEN_259; // @[lut_mem_online.scala 247:34]
  wire  _GEN_262 = io_inputBit ? 1'h0 : _GEN_261; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_263 = i == 10'h48 ? _GEN_262 : _GEN_261; // @[lut_mem_online.scala 247:34]
  wire  _GEN_264 = io_inputBit ? 1'h0 : _GEN_263; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_265 = i == 10'h91 ? _GEN_264 : _GEN_263; // @[lut_mem_online.scala 247:34]
  wire  _GEN_266 = ~io_inputBit | _GEN_265; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_267 = i == 10'h10b ? _GEN_266 : _GEN_265; // @[lut_mem_online.scala 247:34]
  wire  _GEN_268 = ~io_inputBit ? 1'h0 : _GEN_267; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_269 = i == 10'h10c ? _GEN_268 : _GEN_267; // @[lut_mem_online.scala 247:34]
  wire  _GEN_270 = ~io_inputBit | _GEN_269; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_271 = i == 10'h10d ? _GEN_270 : _GEN_269; // @[lut_mem_online.scala 247:34]
  wire  _GEN_272 = ~io_inputBit ? 1'h0 : _GEN_271; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_273 = i == 10'h10e ? _GEN_272 : _GEN_271; // @[lut_mem_online.scala 247:34]
  wire  _GEN_274 = ~io_inputBit | _GEN_273; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_275 = i == 10'h10f ? _GEN_274 : _GEN_273; // @[lut_mem_online.scala 247:34]
  wire  _GEN_276 = ~io_inputBit ? 1'h0 : _GEN_275; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_277 = i == 10'h110 ? _GEN_276 : _GEN_275; // @[lut_mem_online.scala 247:34]
  wire  _GEN_278 = ~io_inputBit | _GEN_277; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_279 = i == 10'h111 ? _GEN_278 : _GEN_277; // @[lut_mem_online.scala 247:34]
  wire  _GEN_280 = ~io_inputBit ? 1'h0 : _GEN_279; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_281 = i == 10'h112 ? _GEN_280 : _GEN_279; // @[lut_mem_online.scala 247:34]
  wire  _GEN_282 = ~io_inputBit | _GEN_281; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_283 = i == 10'h113 ? _GEN_282 : _GEN_281; // @[lut_mem_online.scala 247:34]
  wire  _GEN_284 = ~io_inputBit ? 1'h0 : _GEN_283; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_285 = i == 10'h114 ? _GEN_284 : _GEN_283; // @[lut_mem_online.scala 247:34]
  wire  _GEN_286 = ~io_inputBit | _GEN_285; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_287 = i == 10'h115 ? _GEN_286 : _GEN_285; // @[lut_mem_online.scala 247:34]
  wire  _GEN_288 = ~io_inputBit ? 1'h0 : _GEN_287; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_289 = i == 10'h116 ? _GEN_288 : _GEN_287; // @[lut_mem_online.scala 247:34]
  wire  _GEN_290 = ~io_inputBit | _GEN_289; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_291 = i == 10'h117 ? _GEN_290 : _GEN_289; // @[lut_mem_online.scala 247:34]
  wire  _GEN_292 = ~io_inputBit ? 1'h0 : _GEN_291; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_293 = i == 10'h118 ? _GEN_292 : _GEN_291; // @[lut_mem_online.scala 247:34]
  wire  _GEN_294 = ~io_inputBit | _GEN_293; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_295 = i == 10'h119 ? _GEN_294 : _GEN_293; // @[lut_mem_online.scala 247:34]
  wire  _GEN_296 = ~io_inputBit ? 1'h0 : _GEN_295; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_297 = i == 10'h11a ? _GEN_296 : _GEN_295; // @[lut_mem_online.scala 247:34]
  wire  _GEN_298 = ~io_inputBit | _GEN_297; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_299 = i == 10'h11b ? _GEN_298 : _GEN_297; // @[lut_mem_online.scala 247:34]
  wire  _GEN_300 = ~io_inputBit ? 1'h0 : _GEN_299; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_301 = i == 10'h11c ? _GEN_300 : _GEN_299; // @[lut_mem_online.scala 247:34]
  wire  _GEN_302 = ~io_inputBit | _GEN_301; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_303 = i == 10'h11d ? _GEN_302 : _GEN_301; // @[lut_mem_online.scala 247:34]
  wire  _GEN_304 = ~io_inputBit ? 1'h0 : _GEN_303; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_305 = i == 10'h11e ? _GEN_304 : _GEN_303; // @[lut_mem_online.scala 247:34]
  wire  _GEN_306 = ~io_inputBit | _GEN_305; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_307 = i == 10'h11f ? _GEN_306 : _GEN_305; // @[lut_mem_online.scala 247:34]
  wire  _GEN_308 = ~io_inputBit ? 1'h0 : _GEN_307; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_309 = i == 10'h120 ? _GEN_308 : _GEN_307; // @[lut_mem_online.scala 247:34]
  wire  _GEN_310 = ~io_inputBit | _GEN_309; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_311 = i == 10'h121 ? _GEN_310 : _GEN_309; // @[lut_mem_online.scala 247:34]
  wire  _GEN_312 = ~io_inputBit ? 1'h0 : _GEN_311; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_313 = i == 10'h122 ? _GEN_312 : _GEN_311; // @[lut_mem_online.scala 247:34]
  wire  _GEN_314 = ~io_inputBit | _GEN_313; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_315 = i == 10'h123 ? _GEN_314 : _GEN_313; // @[lut_mem_online.scala 247:34]
  wire  _GEN_316 = ~io_inputBit | _GEN_315; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_317 = i == 10'h218 ? _GEN_316 : _GEN_315; // @[lut_mem_online.scala 247:34]
  wire  _GEN_318 = io_inputBit ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_319 = i == 10'h218 ? _GEN_318 : _GEN_317; // @[lut_mem_online.scala 247:34]
  wire  _GEN_320 = ~io_inputBit ? 1'h0 : _GEN_319; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_321 = i == 10'h21a ? _GEN_320 : _GEN_319; // @[lut_mem_online.scala 247:34]
  wire  _GEN_322 = io_inputBit | _GEN_321; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_323 = i == 10'h21a ? _GEN_322 : _GEN_321; // @[lut_mem_online.scala 247:34]
  wire  _GEN_324 = ~io_inputBit | _GEN_323; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_325 = i == 10'h21c ? _GEN_324 : _GEN_323; // @[lut_mem_online.scala 247:34]
  wire  _GEN_326 = io_inputBit ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_327 = i == 10'h21c ? _GEN_326 : _GEN_325; // @[lut_mem_online.scala 247:34]
  wire  _GEN_328 = ~io_inputBit ? 1'h0 : _GEN_327; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_329 = i == 10'h21e ? _GEN_328 : _GEN_327; // @[lut_mem_online.scala 247:34]
  wire  _GEN_330 = io_inputBit | _GEN_329; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_331 = i == 10'h21e ? _GEN_330 : _GEN_329; // @[lut_mem_online.scala 247:34]
  wire  _GEN_332 = ~io_inputBit | _GEN_331; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_333 = i == 10'h220 ? _GEN_332 : _GEN_331; // @[lut_mem_online.scala 247:34]
  wire  _GEN_334 = io_inputBit ? 1'h0 : _GEN_333; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_335 = i == 10'h220 ? _GEN_334 : _GEN_333; // @[lut_mem_online.scala 247:34]
  wire  _GEN_336 = ~io_inputBit ? 1'h0 : _GEN_335; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_337 = i == 10'h222 ? _GEN_336 : _GEN_335; // @[lut_mem_online.scala 247:34]
  wire  _GEN_338 = io_inputBit | _GEN_337; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_339 = i == 10'h222 ? _GEN_338 : _GEN_337; // @[lut_mem_online.scala 247:34]
  wire  _GEN_340 = ~io_inputBit | _GEN_339; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_341 = i == 10'h224 ? _GEN_340 : _GEN_339; // @[lut_mem_online.scala 247:34]
  wire  _GEN_342 = io_inputBit ? 1'h0 : _GEN_341; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_343 = i == 10'h224 ? _GEN_342 : _GEN_341; // @[lut_mem_online.scala 247:34]
  wire  _GEN_344 = ~io_inputBit ? 1'h0 : _GEN_343; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_345 = i == 10'h226 ? _GEN_344 : _GEN_343; // @[lut_mem_online.scala 247:34]
  wire  _GEN_346 = io_inputBit | _GEN_345; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_347 = i == 10'h226 ? _GEN_346 : _GEN_345; // @[lut_mem_online.scala 247:34]
  wire  _GEN_348 = ~io_inputBit | _GEN_347; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_349 = i == 10'h228 ? _GEN_348 : _GEN_347; // @[lut_mem_online.scala 247:34]
  wire  _GEN_350 = io_inputBit ? 1'h0 : _GEN_349; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_351 = i == 10'h228 ? _GEN_350 : _GEN_349; // @[lut_mem_online.scala 247:34]
  wire  _GEN_352 = ~io_inputBit ? 1'h0 : _GEN_351; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_353 = i == 10'h22a ? _GEN_352 : _GEN_351; // @[lut_mem_online.scala 247:34]
  wire  _GEN_354 = io_inputBit | _GEN_353; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_355 = i == 10'h22a ? _GEN_354 : _GEN_353; // @[lut_mem_online.scala 247:34]
  wire  _GEN_356 = ~io_inputBit | _GEN_355; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_357 = i == 10'h22c ? _GEN_356 : _GEN_355; // @[lut_mem_online.scala 247:34]
  wire  _GEN_358 = io_inputBit ? 1'h0 : _GEN_357; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_359 = i == 10'h22c ? _GEN_358 : _GEN_357; // @[lut_mem_online.scala 247:34]
  wire  _GEN_360 = ~io_inputBit ? 1'h0 : _GEN_359; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_361 = i == 10'h22e ? _GEN_360 : _GEN_359; // @[lut_mem_online.scala 247:34]
  wire  _GEN_362 = io_inputBit | _GEN_361; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_363 = i == 10'h22e ? _GEN_362 : _GEN_361; // @[lut_mem_online.scala 247:34]
  wire  _GEN_364 = ~io_inputBit | _GEN_363; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_365 = i == 10'h230 ? _GEN_364 : _GEN_363; // @[lut_mem_online.scala 247:34]
  wire  _GEN_366 = io_inputBit ? 1'h0 : _GEN_365; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_367 = i == 10'h230 ? _GEN_366 : _GEN_365; // @[lut_mem_online.scala 247:34]
  wire  _GEN_368 = ~io_inputBit ? 1'h0 : _GEN_367; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_369 = i == 10'h232 ? _GEN_368 : _GEN_367; // @[lut_mem_online.scala 247:34]
  wire  _GEN_370 = io_inputBit | _GEN_369; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_371 = i == 10'h232 ? _GEN_370 : _GEN_369; // @[lut_mem_online.scala 247:34]
  wire  _GEN_372 = ~io_inputBit | _GEN_371; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_373 = i == 10'h234 ? _GEN_372 : _GEN_371; // @[lut_mem_online.scala 247:34]
  wire  _GEN_374 = io_inputBit ? 1'h0 : _GEN_373; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_375 = i == 10'h234 ? _GEN_374 : _GEN_373; // @[lut_mem_online.scala 247:34]
  wire  _GEN_376 = ~io_inputBit ? 1'h0 : _GEN_375; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_377 = i == 10'h236 ? _GEN_376 : _GEN_375; // @[lut_mem_online.scala 247:34]
  wire  _GEN_378 = io_inputBit | _GEN_377; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_379 = i == 10'h236 ? _GEN_378 : _GEN_377; // @[lut_mem_online.scala 247:34]
  wire  _GEN_380 = ~io_inputBit | _GEN_379; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_381 = i == 10'h238 ? _GEN_380 : _GEN_379; // @[lut_mem_online.scala 247:34]
  wire  _GEN_382 = io_inputBit ? 1'h0 : _GEN_381; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_383 = i == 10'h238 ? _GEN_382 : _GEN_381; // @[lut_mem_online.scala 247:34]
  wire  _GEN_384 = ~io_inputBit ? 1'h0 : _GEN_383; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_385 = i == 10'h23a ? _GEN_384 : _GEN_383; // @[lut_mem_online.scala 247:34]
  wire  _GEN_386 = io_inputBit | _GEN_385; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_387 = i == 10'h23a ? _GEN_386 : _GEN_385; // @[lut_mem_online.scala 247:34]
  wire  _GEN_388 = ~io_inputBit | _GEN_387; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_389 = i == 10'h23c ? _GEN_388 : _GEN_387; // @[lut_mem_online.scala 247:34]
  wire  _GEN_390 = io_inputBit ? 1'h0 : _GEN_389; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_391 = i == 10'h23c ? _GEN_390 : _GEN_389; // @[lut_mem_online.scala 247:34]
  wire  _GEN_392 = ~io_inputBit ? 1'h0 : _GEN_391; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_393 = i == 10'h23e ? _GEN_392 : _GEN_391; // @[lut_mem_online.scala 247:34]
  wire  _GEN_394 = io_inputBit | _GEN_393; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_395 = i == 10'h23e ? _GEN_394 : _GEN_393; // @[lut_mem_online.scala 247:34]
  wire  _GEN_396 = ~io_inputBit | _GEN_395; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_397 = i == 10'h240 ? _GEN_396 : _GEN_395; // @[lut_mem_online.scala 247:34]
  wire  _GEN_398 = io_inputBit ? 1'h0 : _GEN_397; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_399 = i == 10'h240 ? _GEN_398 : _GEN_397; // @[lut_mem_online.scala 247:34]
  wire  _GEN_400 = ~io_inputBit ? 1'h0 : _GEN_399; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_401 = i == 10'h242 ? _GEN_400 : _GEN_399; // @[lut_mem_online.scala 247:34]
  wire  _GEN_402 = io_inputBit | _GEN_401; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_403 = i == 10'h242 ? _GEN_402 : _GEN_401; // @[lut_mem_online.scala 247:34]
  wire  _GEN_404 = ~io_inputBit | _GEN_403; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_405 = i == 10'h244 ? _GEN_404 : _GEN_403; // @[lut_mem_online.scala 247:34]
  wire  _GEN_406 = io_inputBit ? 1'h0 : _GEN_405; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_407 = i == 10'h244 ? _GEN_406 : _GEN_405; // @[lut_mem_online.scala 247:34]
  wire  _GEN_408 = ~io_inputBit ? 1'h0 : _GEN_407; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_409 = i == 10'h246 ? _GEN_408 : _GEN_407; // @[lut_mem_online.scala 247:34]
  wire  _GEN_410 = io_inputBit | _GEN_409; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_411 = i == 10'h246 ? _GEN_410 : _GEN_409; // @[lut_mem_online.scala 247:34]
  wire  _GEN_412 = ~io_inputBit | _GEN_411; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_413 = i == 10'h248 ? _GEN_412 : _GEN_411; // @[lut_mem_online.scala 247:34]
  wire  _GEN_414 = io_inputBit ? 1'h0 : _GEN_413; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_415 = i == 10'h248 ? _GEN_414 : _GEN_413; // @[lut_mem_online.scala 247:34]
  wire  _GEN_416 = io_inputBit ? 1'h0 : buffer_5; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_417 = i == 10'h0 ? _GEN_416 : buffer_5; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_418 = io_inputBit ? 1'h0 : _GEN_417; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_419 = i == 10'h1 ? _GEN_418 : _GEN_417; // @[lut_mem_online.scala 247:34]
  wire  _GEN_420 = io_inputBit ? 1'h0 : _GEN_419; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_421 = i == 10'h8 ? _GEN_420 : _GEN_419; // @[lut_mem_online.scala 247:34]
  wire  _GEN_422 = ~io_inputBit ? 1'h0 : _GEN_421; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_423 = i == 10'hf ? _GEN_422 : _GEN_421; // @[lut_mem_online.scala 247:34]
  wire  _GEN_424 = io_inputBit ? 1'h0 : _GEN_423; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_425 = i == 10'h11 ? _GEN_424 : _GEN_423; // @[lut_mem_online.scala 247:34]
  wire  _GEN_426 = ~io_inputBit ? 1'h0 : _GEN_425; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_427 = i == 10'h20 ? _GEN_426 : _GEN_425; // @[lut_mem_online.scala 247:34]
  wire  _GEN_428 = io_inputBit ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_429 = i == 10'h48 ? _GEN_428 : _GEN_427; // @[lut_mem_online.scala 247:34]
  wire  _GEN_430 = ~io_inputBit ? 1'h0 : _GEN_429; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_431 = i == 10'h10b ? _GEN_430 : _GEN_429; // @[lut_mem_online.scala 247:34]
  wire  _GEN_432 = io_inputBit ? 1'h0 : _GEN_431; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_433 = i == 10'h124 ? _GEN_432 : _GEN_431; // @[lut_mem_online.scala 247:34]
  wire  _GEN_434 = ~io_inputBit ? 1'h0 : _GEN_433; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_435 = i == 10'h218 ? _GEN_434 : _GEN_433; // @[lut_mem_online.scala 247:34]
  wire  _GEN_436 = io_inputBit | _GEN_435; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_437 = i == 10'h218 ? _GEN_436 : _GEN_435; // @[lut_mem_online.scala 247:34]
  wire  _GEN_438 = ~io_inputBit | _GEN_437; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_439 = i == 10'h219 ? _GEN_438 : _GEN_437; // @[lut_mem_online.scala 247:34]
  wire  _GEN_440 = io_inputBit ? 1'h0 : _GEN_439; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_441 = i == 10'h219 ? _GEN_440 : _GEN_439; // @[lut_mem_online.scala 247:34]
  wire  _GEN_442 = ~io_inputBit ? 1'h0 : _GEN_441; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_443 = i == 10'h21a ? _GEN_442 : _GEN_441; // @[lut_mem_online.scala 247:34]
  wire  _GEN_444 = io_inputBit | _GEN_443; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_445 = i == 10'h21a ? _GEN_444 : _GEN_443; // @[lut_mem_online.scala 247:34]
  wire  _GEN_446 = ~io_inputBit | _GEN_445; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_447 = i == 10'h21b ? _GEN_446 : _GEN_445; // @[lut_mem_online.scala 247:34]
  wire  _GEN_448 = io_inputBit ? 1'h0 : _GEN_447; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_449 = i == 10'h21b ? _GEN_448 : _GEN_447; // @[lut_mem_online.scala 247:34]
  wire  _GEN_450 = ~io_inputBit ? 1'h0 : _GEN_449; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_451 = i == 10'h21c ? _GEN_450 : _GEN_449; // @[lut_mem_online.scala 247:34]
  wire  _GEN_452 = io_inputBit | _GEN_451; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_453 = i == 10'h21c ? _GEN_452 : _GEN_451; // @[lut_mem_online.scala 247:34]
  wire  _GEN_454 = ~io_inputBit | _GEN_453; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_455 = i == 10'h21d ? _GEN_454 : _GEN_453; // @[lut_mem_online.scala 247:34]
  wire  _GEN_456 = io_inputBit ? 1'h0 : _GEN_455; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_457 = i == 10'h21d ? _GEN_456 : _GEN_455; // @[lut_mem_online.scala 247:34]
  wire  _GEN_458 = ~io_inputBit ? 1'h0 : _GEN_457; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_459 = i == 10'h21e ? _GEN_458 : _GEN_457; // @[lut_mem_online.scala 247:34]
  wire  _GEN_460 = io_inputBit | _GEN_459; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_461 = i == 10'h21e ? _GEN_460 : _GEN_459; // @[lut_mem_online.scala 247:34]
  wire  _GEN_462 = ~io_inputBit | _GEN_461; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_463 = i == 10'h21f ? _GEN_462 : _GEN_461; // @[lut_mem_online.scala 247:34]
  wire  _GEN_464 = io_inputBit ? 1'h0 : _GEN_463; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_465 = i == 10'h21f ? _GEN_464 : _GEN_463; // @[lut_mem_online.scala 247:34]
  wire  _GEN_466 = ~io_inputBit ? 1'h0 : _GEN_465; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_467 = i == 10'h220 ? _GEN_466 : _GEN_465; // @[lut_mem_online.scala 247:34]
  wire  _GEN_468 = io_inputBit | _GEN_467; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_469 = i == 10'h220 ? _GEN_468 : _GEN_467; // @[lut_mem_online.scala 247:34]
  wire  _GEN_470 = ~io_inputBit | _GEN_469; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_471 = i == 10'h221 ? _GEN_470 : _GEN_469; // @[lut_mem_online.scala 247:34]
  wire  _GEN_472 = io_inputBit ? 1'h0 : _GEN_471; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_473 = i == 10'h221 ? _GEN_472 : _GEN_471; // @[lut_mem_online.scala 247:34]
  wire  _GEN_474 = ~io_inputBit ? 1'h0 : _GEN_473; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_475 = i == 10'h222 ? _GEN_474 : _GEN_473; // @[lut_mem_online.scala 247:34]
  wire  _GEN_476 = io_inputBit | _GEN_475; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_477 = i == 10'h222 ? _GEN_476 : _GEN_475; // @[lut_mem_online.scala 247:34]
  wire  _GEN_478 = ~io_inputBit | _GEN_477; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_479 = i == 10'h223 ? _GEN_478 : _GEN_477; // @[lut_mem_online.scala 247:34]
  wire  _GEN_480 = io_inputBit ? 1'h0 : _GEN_479; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_481 = i == 10'h223 ? _GEN_480 : _GEN_479; // @[lut_mem_online.scala 247:34]
  wire  _GEN_482 = ~io_inputBit ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_483 = i == 10'h224 ? _GEN_482 : _GEN_481; // @[lut_mem_online.scala 247:34]
  wire  _GEN_484 = io_inputBit | _GEN_483; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_485 = i == 10'h224 ? _GEN_484 : _GEN_483; // @[lut_mem_online.scala 247:34]
  wire  _GEN_486 = ~io_inputBit | _GEN_485; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_487 = i == 10'h225 ? _GEN_486 : _GEN_485; // @[lut_mem_online.scala 247:34]
  wire  _GEN_488 = io_inputBit ? 1'h0 : _GEN_487; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_489 = i == 10'h225 ? _GEN_488 : _GEN_487; // @[lut_mem_online.scala 247:34]
  wire  _GEN_490 = ~io_inputBit ? 1'h0 : _GEN_489; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_491 = i == 10'h226 ? _GEN_490 : _GEN_489; // @[lut_mem_online.scala 247:34]
  wire  _GEN_492 = io_inputBit | _GEN_491; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_493 = i == 10'h226 ? _GEN_492 : _GEN_491; // @[lut_mem_online.scala 247:34]
  wire  _GEN_494 = ~io_inputBit | _GEN_493; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_495 = i == 10'h227 ? _GEN_494 : _GEN_493; // @[lut_mem_online.scala 247:34]
  wire  _GEN_496 = io_inputBit ? 1'h0 : _GEN_495; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_497 = i == 10'h227 ? _GEN_496 : _GEN_495; // @[lut_mem_online.scala 247:34]
  wire  _GEN_498 = ~io_inputBit ? 1'h0 : _GEN_497; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_499 = i == 10'h228 ? _GEN_498 : _GEN_497; // @[lut_mem_online.scala 247:34]
  wire  _GEN_500 = io_inputBit | _GEN_499; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_501 = i == 10'h228 ? _GEN_500 : _GEN_499; // @[lut_mem_online.scala 247:34]
  wire  _GEN_502 = ~io_inputBit | _GEN_501; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_503 = i == 10'h229 ? _GEN_502 : _GEN_501; // @[lut_mem_online.scala 247:34]
  wire  _GEN_504 = io_inputBit ? 1'h0 : _GEN_503; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_505 = i == 10'h229 ? _GEN_504 : _GEN_503; // @[lut_mem_online.scala 247:34]
  wire  _GEN_506 = ~io_inputBit ? 1'h0 : _GEN_505; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_507 = i == 10'h22a ? _GEN_506 : _GEN_505; // @[lut_mem_online.scala 247:34]
  wire  _GEN_508 = io_inputBit | _GEN_507; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_509 = i == 10'h22a ? _GEN_508 : _GEN_507; // @[lut_mem_online.scala 247:34]
  wire  _GEN_510 = ~io_inputBit | _GEN_509; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_511 = i == 10'h22b ? _GEN_510 : _GEN_509; // @[lut_mem_online.scala 247:34]
  wire  _GEN_512 = io_inputBit ? 1'h0 : _GEN_511; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_513 = i == 10'h22b ? _GEN_512 : _GEN_511; // @[lut_mem_online.scala 247:34]
  wire  _GEN_514 = ~io_inputBit ? 1'h0 : _GEN_513; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_515 = i == 10'h22c ? _GEN_514 : _GEN_513; // @[lut_mem_online.scala 247:34]
  wire  _GEN_516 = io_inputBit | _GEN_515; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_517 = i == 10'h22c ? _GEN_516 : _GEN_515; // @[lut_mem_online.scala 247:34]
  wire  _GEN_518 = ~io_inputBit | _GEN_517; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_519 = i == 10'h22d ? _GEN_518 : _GEN_517; // @[lut_mem_online.scala 247:34]
  wire  _GEN_520 = io_inputBit ? 1'h0 : _GEN_519; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_521 = i == 10'h22d ? _GEN_520 : _GEN_519; // @[lut_mem_online.scala 247:34]
  wire  _GEN_522 = ~io_inputBit ? 1'h0 : _GEN_521; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_523 = i == 10'h22e ? _GEN_522 : _GEN_521; // @[lut_mem_online.scala 247:34]
  wire  _GEN_524 = io_inputBit | _GEN_523; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_525 = i == 10'h22e ? _GEN_524 : _GEN_523; // @[lut_mem_online.scala 247:34]
  wire  _GEN_526 = ~io_inputBit | _GEN_525; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_527 = i == 10'h22f ? _GEN_526 : _GEN_525; // @[lut_mem_online.scala 247:34]
  wire  _GEN_528 = io_inputBit ? 1'h0 : _GEN_527; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_529 = i == 10'h22f ? _GEN_528 : _GEN_527; // @[lut_mem_online.scala 247:34]
  wire  _GEN_530 = ~io_inputBit ? 1'h0 : _GEN_529; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_531 = i == 10'h230 ? _GEN_530 : _GEN_529; // @[lut_mem_online.scala 247:34]
  wire  _GEN_532 = io_inputBit | _GEN_531; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_533 = i == 10'h230 ? _GEN_532 : _GEN_531; // @[lut_mem_online.scala 247:34]
  wire  _GEN_534 = ~io_inputBit | _GEN_533; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_535 = i == 10'h231 ? _GEN_534 : _GEN_533; // @[lut_mem_online.scala 247:34]
  wire  _GEN_536 = io_inputBit ? 1'h0 : _GEN_535; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_537 = i == 10'h231 ? _GEN_536 : _GEN_535; // @[lut_mem_online.scala 247:34]
  wire  _GEN_538 = ~io_inputBit ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_539 = i == 10'h232 ? _GEN_538 : _GEN_537; // @[lut_mem_online.scala 247:34]
  wire  _GEN_540 = io_inputBit | _GEN_539; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_541 = i == 10'h232 ? _GEN_540 : _GEN_539; // @[lut_mem_online.scala 247:34]
  wire  _GEN_542 = ~io_inputBit | _GEN_541; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_543 = i == 10'h233 ? _GEN_542 : _GEN_541; // @[lut_mem_online.scala 247:34]
  wire  _GEN_544 = io_inputBit ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_545 = i == 10'h233 ? _GEN_544 : _GEN_543; // @[lut_mem_online.scala 247:34]
  wire  _GEN_546 = ~io_inputBit ? 1'h0 : _GEN_545; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_547 = i == 10'h234 ? _GEN_546 : _GEN_545; // @[lut_mem_online.scala 247:34]
  wire  _GEN_548 = io_inputBit | _GEN_547; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_549 = i == 10'h234 ? _GEN_548 : _GEN_547; // @[lut_mem_online.scala 247:34]
  wire  _GEN_550 = ~io_inputBit | _GEN_549; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_551 = i == 10'h235 ? _GEN_550 : _GEN_549; // @[lut_mem_online.scala 247:34]
  wire  _GEN_552 = io_inputBit ? 1'h0 : _GEN_551; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_553 = i == 10'h235 ? _GEN_552 : _GEN_551; // @[lut_mem_online.scala 247:34]
  wire  _GEN_554 = ~io_inputBit ? 1'h0 : _GEN_553; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_555 = i == 10'h236 ? _GEN_554 : _GEN_553; // @[lut_mem_online.scala 247:34]
  wire  _GEN_556 = io_inputBit | _GEN_555; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_557 = i == 10'h236 ? _GEN_556 : _GEN_555; // @[lut_mem_online.scala 247:34]
  wire  _GEN_558 = ~io_inputBit | _GEN_557; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_559 = i == 10'h237 ? _GEN_558 : _GEN_557; // @[lut_mem_online.scala 247:34]
  wire  _GEN_560 = io_inputBit ? 1'h0 : _GEN_559; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_561 = i == 10'h237 ? _GEN_560 : _GEN_559; // @[lut_mem_online.scala 247:34]
  wire  _GEN_562 = ~io_inputBit ? 1'h0 : _GEN_561; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_563 = i == 10'h238 ? _GEN_562 : _GEN_561; // @[lut_mem_online.scala 247:34]
  wire  _GEN_564 = io_inputBit | _GEN_563; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_565 = i == 10'h238 ? _GEN_564 : _GEN_563; // @[lut_mem_online.scala 247:34]
  wire  _GEN_566 = ~io_inputBit | _GEN_565; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_567 = i == 10'h239 ? _GEN_566 : _GEN_565; // @[lut_mem_online.scala 247:34]
  wire  _GEN_568 = io_inputBit ? 1'h0 : _GEN_567; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_569 = i == 10'h239 ? _GEN_568 : _GEN_567; // @[lut_mem_online.scala 247:34]
  wire  _GEN_570 = ~io_inputBit ? 1'h0 : _GEN_569; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_571 = i == 10'h23a ? _GEN_570 : _GEN_569; // @[lut_mem_online.scala 247:34]
  wire  _GEN_572 = io_inputBit | _GEN_571; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_573 = i == 10'h23a ? _GEN_572 : _GEN_571; // @[lut_mem_online.scala 247:34]
  wire  _GEN_574 = ~io_inputBit | _GEN_573; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_575 = i == 10'h23b ? _GEN_574 : _GEN_573; // @[lut_mem_online.scala 247:34]
  wire  _GEN_576 = io_inputBit ? 1'h0 : _GEN_575; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_577 = i == 10'h23b ? _GEN_576 : _GEN_575; // @[lut_mem_online.scala 247:34]
  wire  _GEN_578 = ~io_inputBit ? 1'h0 : _GEN_577; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_579 = i == 10'h23c ? _GEN_578 : _GEN_577; // @[lut_mem_online.scala 247:34]
  wire  _GEN_580 = io_inputBit | _GEN_579; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_581 = i == 10'h23c ? _GEN_580 : _GEN_579; // @[lut_mem_online.scala 247:34]
  wire  _GEN_582 = ~io_inputBit | _GEN_581; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_583 = i == 10'h23d ? _GEN_582 : _GEN_581; // @[lut_mem_online.scala 247:34]
  wire  _GEN_584 = io_inputBit ? 1'h0 : _GEN_583; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_585 = i == 10'h23d ? _GEN_584 : _GEN_583; // @[lut_mem_online.scala 247:34]
  wire  _GEN_586 = ~io_inputBit ? 1'h0 : _GEN_585; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_587 = i == 10'h23e ? _GEN_586 : _GEN_585; // @[lut_mem_online.scala 247:34]
  wire  _GEN_588 = io_inputBit | _GEN_587; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_589 = i == 10'h23e ? _GEN_588 : _GEN_587; // @[lut_mem_online.scala 247:34]
  wire  _GEN_590 = ~io_inputBit | _GEN_589; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_591 = i == 10'h23f ? _GEN_590 : _GEN_589; // @[lut_mem_online.scala 247:34]
  wire  _GEN_592 = io_inputBit ? 1'h0 : _GEN_591; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_593 = i == 10'h23f ? _GEN_592 : _GEN_591; // @[lut_mem_online.scala 247:34]
  wire  _GEN_594 = ~io_inputBit ? 1'h0 : _GEN_593; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_595 = i == 10'h240 ? _GEN_594 : _GEN_593; // @[lut_mem_online.scala 247:34]
  wire  _GEN_596 = io_inputBit | _GEN_595; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_597 = i == 10'h240 ? _GEN_596 : _GEN_595; // @[lut_mem_online.scala 247:34]
  wire  _GEN_598 = ~io_inputBit | _GEN_597; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_599 = i == 10'h241 ? _GEN_598 : _GEN_597; // @[lut_mem_online.scala 247:34]
  wire  _GEN_600 = io_inputBit ? 1'h0 : _GEN_599; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_601 = i == 10'h241 ? _GEN_600 : _GEN_599; // @[lut_mem_online.scala 247:34]
  wire  _GEN_602 = ~io_inputBit ? 1'h0 : _GEN_601; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_603 = i == 10'h242 ? _GEN_602 : _GEN_601; // @[lut_mem_online.scala 247:34]
  wire  _GEN_604 = io_inputBit | _GEN_603; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_605 = i == 10'h242 ? _GEN_604 : _GEN_603; // @[lut_mem_online.scala 247:34]
  wire  _GEN_606 = ~io_inputBit | _GEN_605; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_607 = i == 10'h243 ? _GEN_606 : _GEN_605; // @[lut_mem_online.scala 247:34]
  wire  _GEN_608 = io_inputBit ? 1'h0 : _GEN_607; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_609 = i == 10'h243 ? _GEN_608 : _GEN_607; // @[lut_mem_online.scala 247:34]
  wire  _GEN_610 = ~io_inputBit ? 1'h0 : _GEN_609; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_611 = i == 10'h244 ? _GEN_610 : _GEN_609; // @[lut_mem_online.scala 247:34]
  wire  _GEN_612 = io_inputBit | _GEN_611; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_613 = i == 10'h244 ? _GEN_612 : _GEN_611; // @[lut_mem_online.scala 247:34]
  wire  _GEN_614 = ~io_inputBit | _GEN_613; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_615 = i == 10'h245 ? _GEN_614 : _GEN_613; // @[lut_mem_online.scala 247:34]
  wire  _GEN_616 = io_inputBit ? 1'h0 : _GEN_615; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_617 = i == 10'h245 ? _GEN_616 : _GEN_615; // @[lut_mem_online.scala 247:34]
  wire  _GEN_618 = ~io_inputBit ? 1'h0 : _GEN_617; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_619 = i == 10'h246 ? _GEN_618 : _GEN_617; // @[lut_mem_online.scala 247:34]
  wire  _GEN_620 = io_inputBit | _GEN_619; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_621 = i == 10'h246 ? _GEN_620 : _GEN_619; // @[lut_mem_online.scala 247:34]
  wire  _GEN_622 = ~io_inputBit | _GEN_621; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_623 = i == 10'h247 ? _GEN_622 : _GEN_621; // @[lut_mem_online.scala 247:34]
  wire  _GEN_624 = io_inputBit ? 1'h0 : _GEN_623; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_625 = i == 10'h247 ? _GEN_624 : _GEN_623; // @[lut_mem_online.scala 247:34]
  wire  _GEN_626 = ~io_inputBit ? 1'h0 : _GEN_625; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_627 = i == 10'h248 ? _GEN_626 : _GEN_625; // @[lut_mem_online.scala 247:34]
  wire  _GEN_628 = io_inputBit | _GEN_627; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_629 = i == 10'h248 ? _GEN_628 : _GEN_627; // @[lut_mem_online.scala 247:34]
  wire  _GEN_630 = ~io_inputBit | _GEN_629; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_631 = i == 10'h249 ? _GEN_630 : _GEN_629; // @[lut_mem_online.scala 247:34]
  wire  _GEN_632 = io_inputBit ? 1'h0 : _GEN_631; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_633 = i == 10'h249 ? _GEN_632 : _GEN_631; // @[lut_mem_online.scala 247:34]
  wire  _GEN_634 = io_inputBit ? 1'h0 : buffer_6; // @[lut_mem_online.scala 219:19 249:46 251:32]
  wire  _GEN_635 = i == 10'h0 ? _GEN_634 : buffer_6; // @[lut_mem_online.scala 219:19 247:34]
  wire  _GEN_636 = io_inputBit ? 1'h0 : _GEN_635; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_637 = i == 10'h1 ? _GEN_636 : _GEN_635; // @[lut_mem_online.scala 247:34]
  wire  _GEN_638 = io_inputBit ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_639 = i == 10'h8 ? _GEN_638 : _GEN_637; // @[lut_mem_online.scala 247:34]
  wire  _GEN_640 = ~io_inputBit ? 1'h0 : _GEN_639; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_641 = i == 10'hf ? _GEN_640 : _GEN_639; // @[lut_mem_online.scala 247:34]
  wire  _GEN_642 = io_inputBit ? 1'h0 : _GEN_641; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_643 = i == 10'h11 ? _GEN_642 : _GEN_641; // @[lut_mem_online.scala 247:34]
  wire  _GEN_644 = ~io_inputBit ? 1'h0 : _GEN_643; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_645 = i == 10'h20 ? _GEN_644 : _GEN_643; // @[lut_mem_online.scala 247:34]
  wire  _GEN_646 = io_inputBit ? 1'h0 : _GEN_645; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_647 = i == 10'h48 ? _GEN_646 : _GEN_645; // @[lut_mem_online.scala 247:34]
  wire  _GEN_648 = ~io_inputBit ? 1'h0 : _GEN_647; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_649 = i == 10'h10b ? _GEN_648 : _GEN_647; // @[lut_mem_online.scala 247:34]
  wire  _GEN_650 = io_inputBit ? 1'h0 : _GEN_649; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_651 = i == 10'h124 ? _GEN_650 : _GEN_649; // @[lut_mem_online.scala 247:34]
  wire  _GEN_652 = ~io_inputBit ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_653 = i == 10'h218 ? _GEN_652 : _GEN_651; // @[lut_mem_online.scala 247:34]
  wire  _GEN_654 = io_inputBit | _GEN_653; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_655 = i == 10'h218 ? _GEN_654 : _GEN_653; // @[lut_mem_online.scala 247:34]
  wire  _GEN_656 = ~io_inputBit ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_657 = i == 10'h219 ? _GEN_656 : _GEN_655; // @[lut_mem_online.scala 247:34]
  wire  _GEN_658 = io_inputBit | _GEN_657; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_659 = i == 10'h219 ? _GEN_658 : _GEN_657; // @[lut_mem_online.scala 247:34]
  wire  _GEN_660 = ~io_inputBit ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_661 = i == 10'h21a ? _GEN_660 : _GEN_659; // @[lut_mem_online.scala 247:34]
  wire  _GEN_662 = io_inputBit | _GEN_661; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_663 = i == 10'h21a ? _GEN_662 : _GEN_661; // @[lut_mem_online.scala 247:34]
  wire  _GEN_664 = ~io_inputBit ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_665 = i == 10'h21b ? _GEN_664 : _GEN_663; // @[lut_mem_online.scala 247:34]
  wire  _GEN_666 = io_inputBit | _GEN_665; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_667 = i == 10'h21b ? _GEN_666 : _GEN_665; // @[lut_mem_online.scala 247:34]
  wire  _GEN_668 = ~io_inputBit ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_669 = i == 10'h21c ? _GEN_668 : _GEN_667; // @[lut_mem_online.scala 247:34]
  wire  _GEN_670 = io_inputBit | _GEN_669; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_671 = i == 10'h21c ? _GEN_670 : _GEN_669; // @[lut_mem_online.scala 247:34]
  wire  _GEN_672 = ~io_inputBit ? 1'h0 : _GEN_671; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_673 = i == 10'h21d ? _GEN_672 : _GEN_671; // @[lut_mem_online.scala 247:34]
  wire  _GEN_674 = io_inputBit | _GEN_673; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_675 = i == 10'h21d ? _GEN_674 : _GEN_673; // @[lut_mem_online.scala 247:34]
  wire  _GEN_676 = ~io_inputBit ? 1'h0 : _GEN_675; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_677 = i == 10'h21e ? _GEN_676 : _GEN_675; // @[lut_mem_online.scala 247:34]
  wire  _GEN_678 = io_inputBit | _GEN_677; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_679 = i == 10'h21e ? _GEN_678 : _GEN_677; // @[lut_mem_online.scala 247:34]
  wire  _GEN_680 = ~io_inputBit ? 1'h0 : _GEN_679; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_681 = i == 10'h21f ? _GEN_680 : _GEN_679; // @[lut_mem_online.scala 247:34]
  wire  _GEN_682 = io_inputBit | _GEN_681; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_683 = i == 10'h21f ? _GEN_682 : _GEN_681; // @[lut_mem_online.scala 247:34]
  wire  _GEN_684 = ~io_inputBit ? 1'h0 : _GEN_683; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_685 = i == 10'h220 ? _GEN_684 : _GEN_683; // @[lut_mem_online.scala 247:34]
  wire  _GEN_686 = io_inputBit | _GEN_685; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_687 = i == 10'h220 ? _GEN_686 : _GEN_685; // @[lut_mem_online.scala 247:34]
  wire  _GEN_688 = ~io_inputBit ? 1'h0 : _GEN_687; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_689 = i == 10'h221 ? _GEN_688 : _GEN_687; // @[lut_mem_online.scala 247:34]
  wire  _GEN_690 = io_inputBit | _GEN_689; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_691 = i == 10'h221 ? _GEN_690 : _GEN_689; // @[lut_mem_online.scala 247:34]
  wire  _GEN_692 = ~io_inputBit ? 1'h0 : _GEN_691; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_693 = i == 10'h222 ? _GEN_692 : _GEN_691; // @[lut_mem_online.scala 247:34]
  wire  _GEN_694 = io_inputBit | _GEN_693; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_695 = i == 10'h222 ? _GEN_694 : _GEN_693; // @[lut_mem_online.scala 247:34]
  wire  _GEN_696 = ~io_inputBit ? 1'h0 : _GEN_695; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_697 = i == 10'h223 ? _GEN_696 : _GEN_695; // @[lut_mem_online.scala 247:34]
  wire  _GEN_698 = io_inputBit | _GEN_697; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_699 = i == 10'h223 ? _GEN_698 : _GEN_697; // @[lut_mem_online.scala 247:34]
  wire  _GEN_700 = ~io_inputBit ? 1'h0 : _GEN_699; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_701 = i == 10'h224 ? _GEN_700 : _GEN_699; // @[lut_mem_online.scala 247:34]
  wire  _GEN_702 = io_inputBit | _GEN_701; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_703 = i == 10'h224 ? _GEN_702 : _GEN_701; // @[lut_mem_online.scala 247:34]
  wire  _GEN_704 = ~io_inputBit ? 1'h0 : _GEN_703; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_705 = i == 10'h225 ? _GEN_704 : _GEN_703; // @[lut_mem_online.scala 247:34]
  wire  _GEN_706 = io_inputBit | _GEN_705; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_707 = i == 10'h225 ? _GEN_706 : _GEN_705; // @[lut_mem_online.scala 247:34]
  wire  _GEN_708 = ~io_inputBit ? 1'h0 : _GEN_707; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_709 = i == 10'h226 ? _GEN_708 : _GEN_707; // @[lut_mem_online.scala 247:34]
  wire  _GEN_710 = io_inputBit | _GEN_709; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_711 = i == 10'h226 ? _GEN_710 : _GEN_709; // @[lut_mem_online.scala 247:34]
  wire  _GEN_712 = ~io_inputBit ? 1'h0 : _GEN_711; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_713 = i == 10'h227 ? _GEN_712 : _GEN_711; // @[lut_mem_online.scala 247:34]
  wire  _GEN_714 = io_inputBit | _GEN_713; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_715 = i == 10'h227 ? _GEN_714 : _GEN_713; // @[lut_mem_online.scala 247:34]
  wire  _GEN_716 = ~io_inputBit ? 1'h0 : _GEN_715; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_717 = i == 10'h228 ? _GEN_716 : _GEN_715; // @[lut_mem_online.scala 247:34]
  wire  _GEN_718 = io_inputBit | _GEN_717; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_719 = i == 10'h228 ? _GEN_718 : _GEN_717; // @[lut_mem_online.scala 247:34]
  wire  _GEN_720 = ~io_inputBit ? 1'h0 : _GEN_719; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_721 = i == 10'h229 ? _GEN_720 : _GEN_719; // @[lut_mem_online.scala 247:34]
  wire  _GEN_722 = io_inputBit | _GEN_721; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_723 = i == 10'h229 ? _GEN_722 : _GEN_721; // @[lut_mem_online.scala 247:34]
  wire  _GEN_724 = ~io_inputBit ? 1'h0 : _GEN_723; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_725 = i == 10'h22a ? _GEN_724 : _GEN_723; // @[lut_mem_online.scala 247:34]
  wire  _GEN_726 = io_inputBit | _GEN_725; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_727 = i == 10'h22a ? _GEN_726 : _GEN_725; // @[lut_mem_online.scala 247:34]
  wire  _GEN_728 = ~io_inputBit ? 1'h0 : _GEN_727; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_729 = i == 10'h22b ? _GEN_728 : _GEN_727; // @[lut_mem_online.scala 247:34]
  wire  _GEN_730 = io_inputBit | _GEN_729; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_731 = i == 10'h22b ? _GEN_730 : _GEN_729; // @[lut_mem_online.scala 247:34]
  wire  _GEN_732 = ~io_inputBit ? 1'h0 : _GEN_731; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_733 = i == 10'h22c ? _GEN_732 : _GEN_731; // @[lut_mem_online.scala 247:34]
  wire  _GEN_734 = io_inputBit | _GEN_733; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_735 = i == 10'h22c ? _GEN_734 : _GEN_733; // @[lut_mem_online.scala 247:34]
  wire  _GEN_736 = ~io_inputBit ? 1'h0 : _GEN_735; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_737 = i == 10'h22d ? _GEN_736 : _GEN_735; // @[lut_mem_online.scala 247:34]
  wire  _GEN_738 = io_inputBit | _GEN_737; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_739 = i == 10'h22d ? _GEN_738 : _GEN_737; // @[lut_mem_online.scala 247:34]
  wire  _GEN_740 = ~io_inputBit ? 1'h0 : _GEN_739; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_741 = i == 10'h22e ? _GEN_740 : _GEN_739; // @[lut_mem_online.scala 247:34]
  wire  _GEN_742 = io_inputBit | _GEN_741; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_743 = i == 10'h22e ? _GEN_742 : _GEN_741; // @[lut_mem_online.scala 247:34]
  wire  _GEN_744 = ~io_inputBit ? 1'h0 : _GEN_743; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_745 = i == 10'h22f ? _GEN_744 : _GEN_743; // @[lut_mem_online.scala 247:34]
  wire  _GEN_746 = io_inputBit | _GEN_745; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_747 = i == 10'h22f ? _GEN_746 : _GEN_745; // @[lut_mem_online.scala 247:34]
  wire  _GEN_748 = ~io_inputBit ? 1'h0 : _GEN_747; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_749 = i == 10'h230 ? _GEN_748 : _GEN_747; // @[lut_mem_online.scala 247:34]
  wire  _GEN_750 = io_inputBit | _GEN_749; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_751 = i == 10'h230 ? _GEN_750 : _GEN_749; // @[lut_mem_online.scala 247:34]
  wire  _GEN_752 = ~io_inputBit ? 1'h0 : _GEN_751; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_753 = i == 10'h231 ? _GEN_752 : _GEN_751; // @[lut_mem_online.scala 247:34]
  wire  _GEN_754 = io_inputBit | _GEN_753; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_755 = i == 10'h231 ? _GEN_754 : _GEN_753; // @[lut_mem_online.scala 247:34]
  wire  _GEN_756 = ~io_inputBit ? 1'h0 : _GEN_755; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_757 = i == 10'h232 ? _GEN_756 : _GEN_755; // @[lut_mem_online.scala 247:34]
  wire  _GEN_758 = io_inputBit | _GEN_757; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_759 = i == 10'h232 ? _GEN_758 : _GEN_757; // @[lut_mem_online.scala 247:34]
  wire  _GEN_760 = ~io_inputBit ? 1'h0 : _GEN_759; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_761 = i == 10'h233 ? _GEN_760 : _GEN_759; // @[lut_mem_online.scala 247:34]
  wire  _GEN_762 = io_inputBit | _GEN_761; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_763 = i == 10'h233 ? _GEN_762 : _GEN_761; // @[lut_mem_online.scala 247:34]
  wire  _GEN_764 = ~io_inputBit ? 1'h0 : _GEN_763; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_765 = i == 10'h234 ? _GEN_764 : _GEN_763; // @[lut_mem_online.scala 247:34]
  wire  _GEN_766 = io_inputBit | _GEN_765; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_767 = i == 10'h234 ? _GEN_766 : _GEN_765; // @[lut_mem_online.scala 247:34]
  wire  _GEN_768 = ~io_inputBit ? 1'h0 : _GEN_767; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_769 = i == 10'h235 ? _GEN_768 : _GEN_767; // @[lut_mem_online.scala 247:34]
  wire  _GEN_770 = io_inputBit | _GEN_769; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_771 = i == 10'h235 ? _GEN_770 : _GEN_769; // @[lut_mem_online.scala 247:34]
  wire  _GEN_772 = ~io_inputBit ? 1'h0 : _GEN_771; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_773 = i == 10'h236 ? _GEN_772 : _GEN_771; // @[lut_mem_online.scala 247:34]
  wire  _GEN_774 = io_inputBit | _GEN_773; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_775 = i == 10'h236 ? _GEN_774 : _GEN_773; // @[lut_mem_online.scala 247:34]
  wire  _GEN_776 = ~io_inputBit ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_777 = i == 10'h237 ? _GEN_776 : _GEN_775; // @[lut_mem_online.scala 247:34]
  wire  _GEN_778 = io_inputBit | _GEN_777; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_779 = i == 10'h237 ? _GEN_778 : _GEN_777; // @[lut_mem_online.scala 247:34]
  wire  _GEN_780 = ~io_inputBit ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_781 = i == 10'h238 ? _GEN_780 : _GEN_779; // @[lut_mem_online.scala 247:34]
  wire  _GEN_782 = io_inputBit | _GEN_781; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_783 = i == 10'h238 ? _GEN_782 : _GEN_781; // @[lut_mem_online.scala 247:34]
  wire  _GEN_784 = ~io_inputBit ? 1'h0 : _GEN_783; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_785 = i == 10'h239 ? _GEN_784 : _GEN_783; // @[lut_mem_online.scala 247:34]
  wire  _GEN_786 = io_inputBit | _GEN_785; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_787 = i == 10'h239 ? _GEN_786 : _GEN_785; // @[lut_mem_online.scala 247:34]
  wire  _GEN_788 = ~io_inputBit ? 1'h0 : _GEN_787; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_789 = i == 10'h23a ? _GEN_788 : _GEN_787; // @[lut_mem_online.scala 247:34]
  wire  _GEN_790 = io_inputBit | _GEN_789; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_791 = i == 10'h23a ? _GEN_790 : _GEN_789; // @[lut_mem_online.scala 247:34]
  wire  _GEN_792 = ~io_inputBit ? 1'h0 : _GEN_791; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_793 = i == 10'h23b ? _GEN_792 : _GEN_791; // @[lut_mem_online.scala 247:34]
  wire  _GEN_794 = io_inputBit | _GEN_793; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_795 = i == 10'h23b ? _GEN_794 : _GEN_793; // @[lut_mem_online.scala 247:34]
  wire  _GEN_796 = ~io_inputBit ? 1'h0 : _GEN_795; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_797 = i == 10'h23c ? _GEN_796 : _GEN_795; // @[lut_mem_online.scala 247:34]
  wire  _GEN_798 = io_inputBit | _GEN_797; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_799 = i == 10'h23c ? _GEN_798 : _GEN_797; // @[lut_mem_online.scala 247:34]
  wire  _GEN_800 = ~io_inputBit ? 1'h0 : _GEN_799; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_801 = i == 10'h23d ? _GEN_800 : _GEN_799; // @[lut_mem_online.scala 247:34]
  wire  _GEN_802 = io_inputBit | _GEN_801; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_803 = i == 10'h23d ? _GEN_802 : _GEN_801; // @[lut_mem_online.scala 247:34]
  wire  _GEN_804 = ~io_inputBit ? 1'h0 : _GEN_803; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_805 = i == 10'h23e ? _GEN_804 : _GEN_803; // @[lut_mem_online.scala 247:34]
  wire  _GEN_806 = io_inputBit | _GEN_805; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_807 = i == 10'h23e ? _GEN_806 : _GEN_805; // @[lut_mem_online.scala 247:34]
  wire  _GEN_808 = ~io_inputBit ? 1'h0 : _GEN_807; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_809 = i == 10'h23f ? _GEN_808 : _GEN_807; // @[lut_mem_online.scala 247:34]
  wire  _GEN_810 = io_inputBit | _GEN_809; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_811 = i == 10'h23f ? _GEN_810 : _GEN_809; // @[lut_mem_online.scala 247:34]
  wire  _GEN_812 = ~io_inputBit ? 1'h0 : _GEN_811; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_813 = i == 10'h240 ? _GEN_812 : _GEN_811; // @[lut_mem_online.scala 247:34]
  wire  _GEN_814 = io_inputBit | _GEN_813; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_815 = i == 10'h240 ? _GEN_814 : _GEN_813; // @[lut_mem_online.scala 247:34]
  wire  _GEN_816 = ~io_inputBit ? 1'h0 : _GEN_815; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_817 = i == 10'h241 ? _GEN_816 : _GEN_815; // @[lut_mem_online.scala 247:34]
  wire  _GEN_818 = io_inputBit | _GEN_817; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_819 = i == 10'h241 ? _GEN_818 : _GEN_817; // @[lut_mem_online.scala 247:34]
  wire  _GEN_820 = ~io_inputBit ? 1'h0 : _GEN_819; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_821 = i == 10'h242 ? _GEN_820 : _GEN_819; // @[lut_mem_online.scala 247:34]
  wire  _GEN_822 = io_inputBit | _GEN_821; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_823 = i == 10'h242 ? _GEN_822 : _GEN_821; // @[lut_mem_online.scala 247:34]
  wire  _GEN_824 = ~io_inputBit ? 1'h0 : _GEN_823; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_825 = i == 10'h243 ? _GEN_824 : _GEN_823; // @[lut_mem_online.scala 247:34]
  wire  _GEN_826 = io_inputBit | _GEN_825; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_827 = i == 10'h243 ? _GEN_826 : _GEN_825; // @[lut_mem_online.scala 247:34]
  wire  _GEN_828 = ~io_inputBit ? 1'h0 : _GEN_827; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_829 = i == 10'h244 ? _GEN_828 : _GEN_827; // @[lut_mem_online.scala 247:34]
  wire  _GEN_830 = io_inputBit | _GEN_829; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_831 = i == 10'h244 ? _GEN_830 : _GEN_829; // @[lut_mem_online.scala 247:34]
  wire  _GEN_832 = ~io_inputBit ? 1'h0 : _GEN_831; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_833 = i == 10'h245 ? _GEN_832 : _GEN_831; // @[lut_mem_online.scala 247:34]
  wire  _GEN_834 = io_inputBit | _GEN_833; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_835 = i == 10'h245 ? _GEN_834 : _GEN_833; // @[lut_mem_online.scala 247:34]
  wire  _GEN_836 = ~io_inputBit ? 1'h0 : _GEN_835; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_837 = i == 10'h246 ? _GEN_836 : _GEN_835; // @[lut_mem_online.scala 247:34]
  wire  _GEN_838 = io_inputBit | _GEN_837; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_839 = i == 10'h246 ? _GEN_838 : _GEN_837; // @[lut_mem_online.scala 247:34]
  wire  _GEN_840 = ~io_inputBit ? 1'h0 : _GEN_839; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_841 = i == 10'h247 ? _GEN_840 : _GEN_839; // @[lut_mem_online.scala 247:34]
  wire  _GEN_842 = io_inputBit | _GEN_841; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_843 = i == 10'h247 ? _GEN_842 : _GEN_841; // @[lut_mem_online.scala 247:34]
  wire  _GEN_844 = ~io_inputBit ? 1'h0 : _GEN_843; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_845 = i == 10'h248 ? _GEN_844 : _GEN_843; // @[lut_mem_online.scala 247:34]
  wire  _GEN_846 = io_inputBit | _GEN_845; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_847 = i == 10'h248 ? _GEN_846 : _GEN_845; // @[lut_mem_online.scala 247:34]
  wire  _GEN_848 = ~io_inputBit ? 1'h0 : _GEN_847; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_849 = i == 10'h249 ? _GEN_848 : _GEN_847; // @[lut_mem_online.scala 247:34]
  wire  _GEN_850 = io_inputBit | _GEN_849; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_851 = i == 10'h249 ? _GEN_850 : _GEN_849; // @[lut_mem_online.scala 247:34]
  wire  _GEN_852 = io_inputBit ? 1'h0 : _GEN_21; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_853 = i == 10'h0 ? _GEN_852 : _GEN_21; // @[lut_mem_online.scala 247:34]
  wire  _GEN_854 = io_inputBit ? 1'h0 : _GEN_853; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_855 = i == 10'h1 ? _GEN_854 : _GEN_853; // @[lut_mem_online.scala 247:34]
  wire  _GEN_856 = ~io_inputBit ? 1'h0 : _GEN_855; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_857 = i == 10'h7 ? _GEN_856 : _GEN_855; // @[lut_mem_online.scala 247:34]
  wire  _GEN_858 = ~io_inputBit | _GEN_857; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_859 = i == 10'h8 ? _GEN_858 : _GEN_857; // @[lut_mem_online.scala 247:34]
  wire  _GEN_860 = ~io_inputBit ? 1'h0 : _GEN_859; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_861 = i == 10'h10 ? _GEN_860 : _GEN_859; // @[lut_mem_online.scala 247:34]
  wire  _GEN_862 = ~io_inputBit | _GEN_861; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_863 = i == 10'h12 ? _GEN_862 : _GEN_861; // @[lut_mem_online.scala 247:34]
  wire  _GEN_864 = ~io_inputBit ? 1'h0 : _GEN_863; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_865 = i == 10'h22 ? _GEN_864 : _GEN_863; // @[lut_mem_online.scala 247:34]
  wire  _GEN_866 = io_inputBit ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_867 = i == 10'h26 ? _GEN_866 : _GEN_865; // @[lut_mem_online.scala 247:34]
  wire  _GEN_868 = io_inputBit | _GEN_867; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_869 = i == 10'h46 ? _GEN_868 : _GEN_867; // @[lut_mem_online.scala 247:34]
  wire  _GEN_870 = ~io_inputBit | _GEN_869; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_871 = i == 10'h4d ? _GEN_870 : _GEN_869; // @[lut_mem_online.scala 247:34]
  wire  _GEN_872 = io_inputBit | _GEN_871; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_873 = i == 10'h8d ? _GEN_872 : _GEN_871; // @[lut_mem_online.scala 247:34]
  wire  _GEN_874 = ~io_inputBit | _GEN_873; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_875 = i == 10'h9c ? _GEN_874 : _GEN_873; // @[lut_mem_online.scala 247:34]
  wire  _GEN_876 = ~io_inputBit ? 1'h0 : _GEN_875; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_877 = i == 10'h11b ? _GEN_876 : _GEN_875; // @[lut_mem_online.scala 247:34]
  wire  _GEN_878 = io_inputBit | _GEN_877; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_879 = i == 10'h11b ? _GEN_878 : _GEN_877; // @[lut_mem_online.scala 247:34]
  wire  _GEN_880 = io_inputBit ? 1'h0 : _GEN_879; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_881 = i == 10'h13a ? _GEN_880 : _GEN_879; // @[lut_mem_online.scala 247:34]
  wire  _GEN_882 = ~io_inputBit | _GEN_881; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_883 = i == 10'h275 ? _GEN_882 : _GEN_881; // @[lut_mem_online.scala 247:34]
  wire  _GEN_886 = io_inputBit ? 1'h0 : _GEN_65; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_887 = i == 10'h0 ? _GEN_886 : _GEN_65; // @[lut_mem_online.scala 247:34]
  wire  _GEN_888 = io_inputBit ? 1'h0 : _GEN_887; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_889 = i == 10'h4 ? _GEN_888 : _GEN_887; // @[lut_mem_online.scala 247:34]
  wire  _GEN_890 = ~io_inputBit ? 1'h0 : _GEN_889; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_891 = i == 10'h7 ? _GEN_890 : _GEN_889; // @[lut_mem_online.scala 247:34]
  wire  _GEN_892 = io_inputBit ? 1'h0 : _GEN_891; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_893 = i == 10'h9 ? _GEN_892 : _GEN_891; // @[lut_mem_online.scala 247:34]
  wire  _GEN_894 = io_inputBit | _GEN_893; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_895 = i == 10'h11 ? _GEN_894 : _GEN_893; // @[lut_mem_online.scala 247:34]
  wire  _GEN_896 = io_inputBit ? 1'h0 : _GEN_895; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_897 = i == 10'h13 ? _GEN_896 : _GEN_895; // @[lut_mem_online.scala 247:34]
  wire  _GEN_898 = ~io_inputBit ? 1'h0 : _GEN_897; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_899 = i == 10'h21 ? _GEN_898 : _GEN_897; // @[lut_mem_online.scala 247:34]
  wire  _GEN_900 = ~io_inputBit | _GEN_899; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_901 = i == 10'h22 ? _GEN_900 : _GEN_899; // @[lut_mem_online.scala 247:34]
  wire  _GEN_902 = ~io_inputBit ? 1'h0 : _GEN_901; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_903 = i == 10'h23 ? _GEN_902 : _GEN_901; // @[lut_mem_online.scala 247:34]
  wire  _GEN_904 = io_inputBit ? 1'h0 : _GEN_903; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_905 = i == 10'h25 ? _GEN_904 : _GEN_903; // @[lut_mem_online.scala 247:34]
  wire  _GEN_906 = io_inputBit | _GEN_905; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_907 = i == 10'h26 ? _GEN_906 : _GEN_905; // @[lut_mem_online.scala 247:34]
  wire  _GEN_908 = io_inputBit ? 1'h0 : _GEN_907; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_909 = i == 10'h27 ? _GEN_908 : _GEN_907; // @[lut_mem_online.scala 247:34]
  wire  _GEN_910 = io_inputBit | _GEN_909; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_911 = i == 10'h44 ? _GEN_910 : _GEN_909; // @[lut_mem_online.scala 247:34]
  wire  _GEN_912 = io_inputBit ? 1'h0 : _GEN_911; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_913 = i == 10'h46 ? _GEN_912 : _GEN_911; // @[lut_mem_online.scala 247:34]
  wire  _GEN_914 = io_inputBit | _GEN_913; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_915 = i == 10'h48 ? _GEN_914 : _GEN_913; // @[lut_mem_online.scala 247:34]
  wire  _GEN_916 = ~io_inputBit | _GEN_915; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_917 = i == 10'h4b ? _GEN_916 : _GEN_915; // @[lut_mem_online.scala 247:34]
  wire  _GEN_918 = ~io_inputBit ? 1'h0 : _GEN_917; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_919 = i == 10'h4d ? _GEN_918 : _GEN_917; // @[lut_mem_online.scala 247:34]
  wire  _GEN_920 = ~io_inputBit | _GEN_919; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_921 = i == 10'h4f ? _GEN_920 : _GEN_919; // @[lut_mem_online.scala 247:34]
  wire  _GEN_922 = io_inputBit | _GEN_921; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_923 = i == 10'h89 ? _GEN_922 : _GEN_921; // @[lut_mem_online.scala 247:34]
  wire  _GEN_924 = io_inputBit ? 1'h0 : _GEN_923; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_925 = i == 10'h8d ? _GEN_924 : _GEN_923; // @[lut_mem_online.scala 247:34]
  wire  _GEN_926 = io_inputBit | _GEN_925; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_927 = i == 10'h91 ? _GEN_926 : _GEN_925; // @[lut_mem_online.scala 247:34]
  wire  _GEN_928 = ~io_inputBit | _GEN_927; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_929 = i == 10'h98 ? _GEN_928 : _GEN_927; // @[lut_mem_online.scala 247:34]
  wire  _GEN_930 = ~io_inputBit ? 1'h0 : _GEN_929; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_931 = i == 10'h9c ? _GEN_930 : _GEN_929; // @[lut_mem_online.scala 247:34]
  wire  _GEN_932 = ~io_inputBit | _GEN_931; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_933 = i == 10'ha0 ? _GEN_932 : _GEN_931; // @[lut_mem_online.scala 247:34]
  wire  _GEN_934 = ~io_inputBit ? 1'h0 : _GEN_933; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_935 = i == 10'h113 ? _GEN_934 : _GEN_933; // @[lut_mem_online.scala 247:34]
  wire  _GEN_936 = io_inputBit | _GEN_935; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_937 = i == 10'h113 ? _GEN_936 : _GEN_935; // @[lut_mem_online.scala 247:34]
  wire  _GEN_938 = ~io_inputBit | _GEN_937; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_939 = i == 10'h11b ? _GEN_938 : _GEN_937; // @[lut_mem_online.scala 247:34]
  wire  _GEN_940 = io_inputBit ? 1'h0 : _GEN_939; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_941 = i == 10'h11b ? _GEN_940 : _GEN_939; // @[lut_mem_online.scala 247:34]
  wire  _GEN_942 = ~io_inputBit ? 1'h0 : _GEN_941; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_943 = i == 10'h123 ? _GEN_942 : _GEN_941; // @[lut_mem_online.scala 247:34]
  wire  _GEN_944 = io_inputBit | _GEN_943; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_945 = i == 10'h123 ? _GEN_944 : _GEN_943; // @[lut_mem_online.scala 247:34]
  wire  _GEN_946 = io_inputBit ? 1'h0 : _GEN_945; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_947 = i == 10'h132 ? _GEN_946 : _GEN_945; // @[lut_mem_online.scala 247:34]
  wire  _GEN_948 = io_inputBit | _GEN_947; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_949 = i == 10'h13a ? _GEN_948 : _GEN_947; // @[lut_mem_online.scala 247:34]
  wire  _GEN_950 = io_inputBit ? 1'h0 : _GEN_949; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_951 = i == 10'h142 ? _GEN_950 : _GEN_949; // @[lut_mem_online.scala 247:34]
  wire  _GEN_952 = ~io_inputBit | _GEN_951; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_953 = i == 10'h265 ? _GEN_952 : _GEN_951; // @[lut_mem_online.scala 247:34]
  wire  _GEN_954 = io_inputBit ? 1'h0 : _GEN_953; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_955 = i == 10'h265 ? _GEN_954 : _GEN_953; // @[lut_mem_online.scala 247:34]
  wire  _GEN_956 = ~io_inputBit ? 1'h0 : _GEN_955; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_957 = i == 10'h275 ? _GEN_956 : _GEN_955; // @[lut_mem_online.scala 247:34]
  wire  _GEN_958 = io_inputBit | _GEN_957; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_959 = i == 10'h275 ? _GEN_958 : _GEN_957; // @[lut_mem_online.scala 247:34]
  wire  _GEN_960 = ~io_inputBit | _GEN_959; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_961 = i == 10'h285 ? _GEN_960 : _GEN_959; // @[lut_mem_online.scala 247:34]
  wire  _GEN_964 = io_inputBit ? 1'h0 : _GEN_139; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_965 = i == 10'h0 ? _GEN_964 : _GEN_139; // @[lut_mem_online.scala 247:34]
  wire  _GEN_966 = io_inputBit ? 1'h0 : _GEN_965; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_967 = i == 10'h4 ? _GEN_966 : _GEN_965; // @[lut_mem_online.scala 247:34]
  wire  _GEN_968 = ~io_inputBit ? 1'h0 : _GEN_967; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_969 = i == 10'h7 ? _GEN_968 : _GEN_967; // @[lut_mem_online.scala 247:34]
  wire  _GEN_970 = io_inputBit ? 1'h0 : _GEN_969; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_971 = i == 10'h9 ? _GEN_970 : _GEN_969; // @[lut_mem_online.scala 247:34]
  wire  _GEN_972 = io_inputBit ? 1'h0 : _GEN_971; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_973 = i == 10'h11 ? _GEN_972 : _GEN_971; // @[lut_mem_online.scala 247:34]
  wire  _GEN_974 = io_inputBit ? 1'h0 : _GEN_973; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_975 = i == 10'h13 ? _GEN_974 : _GEN_973; // @[lut_mem_online.scala 247:34]
  wire  _GEN_976 = io_inputBit | _GEN_975; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_977 = i == 10'h43 ? _GEN_976 : _GEN_975; // @[lut_mem_online.scala 247:34]
  wire  _GEN_978 = io_inputBit ? 1'h0 : _GEN_977; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_979 = i == 10'h44 ? _GEN_978 : _GEN_977; // @[lut_mem_online.scala 247:34]
  wire  _GEN_980 = io_inputBit | _GEN_979; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_981 = i == 10'h45 ? _GEN_980 : _GEN_979; // @[lut_mem_online.scala 247:34]
  wire  _GEN_982 = io_inputBit ? 1'h0 : _GEN_981; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_983 = i == 10'h46 ? _GEN_982 : _GEN_981; // @[lut_mem_online.scala 247:34]
  wire  _GEN_984 = io_inputBit | _GEN_983; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_985 = i == 10'h47 ? _GEN_984 : _GEN_983; // @[lut_mem_online.scala 247:34]
  wire  _GEN_986 = io_inputBit ? 1'h0 : _GEN_985; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_987 = i == 10'h48 ? _GEN_986 : _GEN_985; // @[lut_mem_online.scala 247:34]
  wire  _GEN_988 = ~io_inputBit ? 1'h0 : _GEN_987; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_989 = i == 10'h4b ? _GEN_988 : _GEN_987; // @[lut_mem_online.scala 247:34]
  wire  _GEN_990 = ~io_inputBit | _GEN_989; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_991 = i == 10'h4c ? _GEN_990 : _GEN_989; // @[lut_mem_online.scala 247:34]
  wire  _GEN_992 = ~io_inputBit ? 1'h0 : _GEN_991; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_993 = i == 10'h4d ? _GEN_992 : _GEN_991; // @[lut_mem_online.scala 247:34]
  wire  _GEN_994 = ~io_inputBit | _GEN_993; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_995 = i == 10'h4e ? _GEN_994 : _GEN_993; // @[lut_mem_online.scala 247:34]
  wire  _GEN_996 = ~io_inputBit ? 1'h0 : _GEN_995; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_997 = i == 10'h4f ? _GEN_996 : _GEN_995; // @[lut_mem_online.scala 247:34]
  wire  _GEN_998 = ~io_inputBit | _GEN_997; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_999 = i == 10'h50 ? _GEN_998 : _GEN_997; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1000 = io_inputBit | _GEN_999; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1001 = i == 10'h87 ? _GEN_1000 : _GEN_999; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1002 = io_inputBit ? 1'h0 : _GEN_1001; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1003 = i == 10'h89 ? _GEN_1002 : _GEN_1001; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1004 = io_inputBit | _GEN_1003; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1005 = i == 10'h8b ? _GEN_1004 : _GEN_1003; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1006 = io_inputBit ? 1'h0 : _GEN_1005; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1007 = i == 10'h8d ? _GEN_1006 : _GEN_1005; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1008 = io_inputBit | _GEN_1007; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1009 = i == 10'h8f ? _GEN_1008 : _GEN_1007; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1010 = io_inputBit ? 1'h0 : _GEN_1009; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1011 = i == 10'h91 ? _GEN_1010 : _GEN_1009; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1012 = ~io_inputBit ? 1'h0 : _GEN_1011; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1013 = i == 10'h98 ? _GEN_1012 : _GEN_1011; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1014 = ~io_inputBit | _GEN_1013; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1015 = i == 10'h9a ? _GEN_1014 : _GEN_1013; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1016 = ~io_inputBit ? 1'h0 : _GEN_1015; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1017 = i == 10'h9c ? _GEN_1016 : _GEN_1015; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1018 = ~io_inputBit | _GEN_1017; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1019 = i == 10'h9e ? _GEN_1018 : _GEN_1017; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1020 = ~io_inputBit ? 1'h0 : _GEN_1019; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1021 = i == 10'ha0 ? _GEN_1020 : _GEN_1019; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1022 = ~io_inputBit | _GEN_1021; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1023 = i == 10'ha2 ? _GEN_1022 : _GEN_1021; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1024 = ~io_inputBit ? 1'h0 : _GEN_1023; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1025 = i == 10'h10f ? _GEN_1024 : _GEN_1023; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1026 = io_inputBit | _GEN_1025; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1027 = i == 10'h10f ? _GEN_1026 : _GEN_1025; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1028 = ~io_inputBit | _GEN_1027; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1029 = i == 10'h113 ? _GEN_1028 : _GEN_1027; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1030 = io_inputBit ? 1'h0 : _GEN_1029; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1031 = i == 10'h113 ? _GEN_1030 : _GEN_1029; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1032 = ~io_inputBit ? 1'h0 : _GEN_1031; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1033 = i == 10'h117 ? _GEN_1032 : _GEN_1031; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1034 = io_inputBit | _GEN_1033; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1035 = i == 10'h117 ? _GEN_1034 : _GEN_1033; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1036 = ~io_inputBit | _GEN_1035; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1037 = i == 10'h11b ? _GEN_1036 : _GEN_1035; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1038 = io_inputBit ? 1'h0 : _GEN_1037; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1039 = i == 10'h11b ? _GEN_1038 : _GEN_1037; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1040 = ~io_inputBit ? 1'h0 : _GEN_1039; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1041 = i == 10'h11f ? _GEN_1040 : _GEN_1039; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1042 = io_inputBit | _GEN_1041; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1043 = i == 10'h11f ? _GEN_1042 : _GEN_1041; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1044 = ~io_inputBit | _GEN_1043; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1045 = i == 10'h123 ? _GEN_1044 : _GEN_1043; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1046 = io_inputBit ? 1'h0 : _GEN_1045; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1047 = i == 10'h123 ? _GEN_1046 : _GEN_1045; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1048 = io_inputBit | _GEN_1047; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1049 = i == 10'h132 ? _GEN_1048 : _GEN_1047; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1050 = io_inputBit ? 1'h0 : _GEN_1049; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1051 = i == 10'h136 ? _GEN_1050 : _GEN_1049; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1052 = io_inputBit | _GEN_1051; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1053 = i == 10'h13a ? _GEN_1052 : _GEN_1051; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1054 = io_inputBit ? 1'h0 : _GEN_1053; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1055 = i == 10'h13e ? _GEN_1054 : _GEN_1053; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1056 = io_inputBit | _GEN_1055; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1057 = i == 10'h142 ? _GEN_1056 : _GEN_1055; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1058 = io_inputBit ? 1'h0 : _GEN_1057; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1059 = i == 10'h146 ? _GEN_1058 : _GEN_1057; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1060 = ~io_inputBit ? 1'h0 : _GEN_1059; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1061 = i == 10'h265 ? _GEN_1060 : _GEN_1059; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1062 = io_inputBit | _GEN_1061; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1063 = i == 10'h265 ? _GEN_1062 : _GEN_1061; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1064 = ~io_inputBit | _GEN_1063; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1065 = i == 10'h26d ? _GEN_1064 : _GEN_1063; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1066 = io_inputBit ? 1'h0 : _GEN_1065; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1067 = i == 10'h26d ? _GEN_1066 : _GEN_1065; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1068 = ~io_inputBit ? 1'h0 : _GEN_1067; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1069 = i == 10'h275 ? _GEN_1068 : _GEN_1067; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1070 = io_inputBit | _GEN_1069; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1071 = i == 10'h275 ? _GEN_1070 : _GEN_1069; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1072 = ~io_inputBit | _GEN_1071; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1073 = i == 10'h27d ? _GEN_1072 : _GEN_1071; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1074 = io_inputBit ? 1'h0 : _GEN_1073; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1075 = i == 10'h27d ? _GEN_1074 : _GEN_1073; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1076 = ~io_inputBit ? 1'h0 : _GEN_1075; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1077 = i == 10'h285 ? _GEN_1076 : _GEN_1075; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1078 = io_inputBit | _GEN_1077; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1079 = i == 10'h285 ? _GEN_1078 : _GEN_1077; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1080 = ~io_inputBit | _GEN_1079; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1081 = i == 10'h28d ? _GEN_1080 : _GEN_1079; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1084 = io_inputBit ? 1'h0 : _GEN_249; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1085 = i == 10'h0 ? _GEN_1084 : _GEN_249; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1086 = io_inputBit ? 1'h0 : _GEN_1085; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1087 = i == 10'h4 ? _GEN_1086 : _GEN_1085; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1088 = io_inputBit ? 1'h0 : _GEN_1087; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1089 = i == 10'h9 ? _GEN_1088 : _GEN_1087; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1090 = ~io_inputBit ? 1'h0 : _GEN_1089; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1091 = i == 10'hf ? _GEN_1090 : _GEN_1089; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1092 = io_inputBit ? 1'h0 : _GEN_1091; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1093 = i == 10'h11 ? _GEN_1092 : _GEN_1091; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1094 = ~io_inputBit ? 1'h0 : _GEN_1093; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1095 = i == 10'h20 ? _GEN_1094 : _GEN_1093; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1096 = io_inputBit ? 1'h0 : _GEN_1095; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1097 = i == 10'h28 ? _GEN_1096 : _GEN_1095; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1098 = ~io_inputBit ? 1'h0 : _GEN_1097; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1099 = i == 10'h42 ? _GEN_1098 : _GEN_1097; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1100 = io_inputBit ? 1'h0 : _GEN_1099; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1101 = i == 10'h48 ? _GEN_1100 : _GEN_1099; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1102 = ~io_inputBit ? 1'h0 : _GEN_1101; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1103 = i == 10'h4b ? _GEN_1102 : _GEN_1101; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1104 = io_inputBit ? 1'h0 : _GEN_1103; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1105 = i == 10'h51 ? _GEN_1104 : _GEN_1103; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1106 = io_inputBit | _GEN_1105; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1107 = i == 10'h86 ? _GEN_1106 : _GEN_1105; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1108 = io_inputBit ? 1'h0 : _GEN_1107; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1109 = i == 10'h87 ? _GEN_1108 : _GEN_1107; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1110 = io_inputBit | _GEN_1109; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1111 = i == 10'h88 ? _GEN_1110 : _GEN_1109; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1112 = io_inputBit ? 1'h0 : _GEN_1111; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1113 = i == 10'h89 ? _GEN_1112 : _GEN_1111; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1114 = io_inputBit | _GEN_1113; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1115 = i == 10'h8a ? _GEN_1114 : _GEN_1113; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1116 = io_inputBit ? 1'h0 : _GEN_1115; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1117 = i == 10'h8b ? _GEN_1116 : _GEN_1115; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1118 = io_inputBit | _GEN_1117; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1119 = i == 10'h8c ? _GEN_1118 : _GEN_1117; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1120 = io_inputBit ? 1'h0 : _GEN_1119; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1121 = i == 10'h8d ? _GEN_1120 : _GEN_1119; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1122 = io_inputBit | _GEN_1121; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1123 = i == 10'h8e ? _GEN_1122 : _GEN_1121; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1124 = io_inputBit ? 1'h0 : _GEN_1123; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1125 = i == 10'h8f ? _GEN_1124 : _GEN_1123; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1126 = io_inputBit | _GEN_1125; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1127 = i == 10'h90 ? _GEN_1126 : _GEN_1125; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1128 = io_inputBit ? 1'h0 : _GEN_1127; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1129 = i == 10'h91 ? _GEN_1128 : _GEN_1127; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1130 = ~io_inputBit ? 1'h0 : _GEN_1129; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1131 = i == 10'h98 ? _GEN_1130 : _GEN_1129; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1132 = ~io_inputBit | _GEN_1131; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1133 = i == 10'h99 ? _GEN_1132 : _GEN_1131; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1134 = ~io_inputBit ? 1'h0 : _GEN_1133; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1135 = i == 10'h9a ? _GEN_1134 : _GEN_1133; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1136 = ~io_inputBit | _GEN_1135; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1137 = i == 10'h9b ? _GEN_1136 : _GEN_1135; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1138 = ~io_inputBit ? 1'h0 : _GEN_1137; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1139 = i == 10'h9c ? _GEN_1138 : _GEN_1137; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1140 = ~io_inputBit | _GEN_1139; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1141 = i == 10'h9d ? _GEN_1140 : _GEN_1139; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1142 = ~io_inputBit ? 1'h0 : _GEN_1141; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1143 = i == 10'h9e ? _GEN_1142 : _GEN_1141; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1144 = ~io_inputBit | _GEN_1143; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1145 = i == 10'h9f ? _GEN_1144 : _GEN_1143; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1146 = ~io_inputBit ? 1'h0 : _GEN_1145; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1147 = i == 10'ha0 ? _GEN_1146 : _GEN_1145; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1148 = ~io_inputBit | _GEN_1147; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1149 = i == 10'ha1 ? _GEN_1148 : _GEN_1147; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1150 = ~io_inputBit ? 1'h0 : _GEN_1149; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1151 = i == 10'ha2 ? _GEN_1150 : _GEN_1149; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1152 = ~io_inputBit | _GEN_1151; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1153 = i == 10'ha3 ? _GEN_1152 : _GEN_1151; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1154 = ~io_inputBit ? 1'h0 : _GEN_1153; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1155 = i == 10'h10d ? _GEN_1154 : _GEN_1153; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1156 = io_inputBit | _GEN_1155; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1157 = i == 10'h10d ? _GEN_1156 : _GEN_1155; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1158 = ~io_inputBit | _GEN_1157; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1159 = i == 10'h10f ? _GEN_1158 : _GEN_1157; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1160 = io_inputBit ? 1'h0 : _GEN_1159; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1161 = i == 10'h10f ? _GEN_1160 : _GEN_1159; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1162 = ~io_inputBit ? 1'h0 : _GEN_1161; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1163 = i == 10'h111 ? _GEN_1162 : _GEN_1161; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1164 = io_inputBit | _GEN_1163; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1165 = i == 10'h111 ? _GEN_1164 : _GEN_1163; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1166 = ~io_inputBit | _GEN_1165; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1167 = i == 10'h113 ? _GEN_1166 : _GEN_1165; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1168 = io_inputBit ? 1'h0 : _GEN_1167; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1169 = i == 10'h113 ? _GEN_1168 : _GEN_1167; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1170 = ~io_inputBit ? 1'h0 : _GEN_1169; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1171 = i == 10'h115 ? _GEN_1170 : _GEN_1169; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1172 = io_inputBit | _GEN_1171; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1173 = i == 10'h115 ? _GEN_1172 : _GEN_1171; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1174 = ~io_inputBit | _GEN_1173; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1175 = i == 10'h117 ? _GEN_1174 : _GEN_1173; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1176 = io_inputBit ? 1'h0 : _GEN_1175; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1177 = i == 10'h117 ? _GEN_1176 : _GEN_1175; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1178 = ~io_inputBit ? 1'h0 : _GEN_1177; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1179 = i == 10'h119 ? _GEN_1178 : _GEN_1177; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1180 = io_inputBit | _GEN_1179; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1181 = i == 10'h119 ? _GEN_1180 : _GEN_1179; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1182 = ~io_inputBit | _GEN_1181; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1183 = i == 10'h11b ? _GEN_1182 : _GEN_1181; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1184 = io_inputBit ? 1'h0 : _GEN_1183; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1185 = i == 10'h11b ? _GEN_1184 : _GEN_1183; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1186 = ~io_inputBit ? 1'h0 : _GEN_1185; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1187 = i == 10'h11d ? _GEN_1186 : _GEN_1185; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1188 = io_inputBit | _GEN_1187; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1189 = i == 10'h11d ? _GEN_1188 : _GEN_1187; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1190 = ~io_inputBit | _GEN_1189; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1191 = i == 10'h11f ? _GEN_1190 : _GEN_1189; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1192 = io_inputBit ? 1'h0 : _GEN_1191; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1193 = i == 10'h11f ? _GEN_1192 : _GEN_1191; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1194 = ~io_inputBit ? 1'h0 : _GEN_1193; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1195 = i == 10'h121 ? _GEN_1194 : _GEN_1193; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1196 = io_inputBit | _GEN_1195; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1197 = i == 10'h121 ? _GEN_1196 : _GEN_1195; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1198 = ~io_inputBit | _GEN_1197; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1199 = i == 10'h123 ? _GEN_1198 : _GEN_1197; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1200 = io_inputBit ? 1'h0 : _GEN_1199; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1201 = i == 10'h123 ? _GEN_1200 : _GEN_1199; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1202 = io_inputBit | _GEN_1201; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1203 = i == 10'h132 ? _GEN_1202 : _GEN_1201; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1204 = io_inputBit ? 1'h0 : _GEN_1203; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1205 = i == 10'h134 ? _GEN_1204 : _GEN_1203; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1206 = io_inputBit | _GEN_1205; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1207 = i == 10'h136 ? _GEN_1206 : _GEN_1205; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1208 = io_inputBit ? 1'h0 : _GEN_1207; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1209 = i == 10'h138 ? _GEN_1208 : _GEN_1207; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1210 = io_inputBit | _GEN_1209; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1211 = i == 10'h13a ? _GEN_1210 : _GEN_1209; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1212 = io_inputBit ? 1'h0 : _GEN_1211; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1213 = i == 10'h13c ? _GEN_1212 : _GEN_1211; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1214 = io_inputBit | _GEN_1213; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1215 = i == 10'h13e ? _GEN_1214 : _GEN_1213; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1216 = io_inputBit ? 1'h0 : _GEN_1215; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1217 = i == 10'h140 ? _GEN_1216 : _GEN_1215; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1218 = io_inputBit | _GEN_1217; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1219 = i == 10'h142 ? _GEN_1218 : _GEN_1217; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1220 = io_inputBit ? 1'h0 : _GEN_1219; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1221 = i == 10'h144 ? _GEN_1220 : _GEN_1219; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1222 = io_inputBit | _GEN_1221; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1223 = i == 10'h146 ? _GEN_1222 : _GEN_1221; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1224 = io_inputBit ? 1'h0 : _GEN_1223; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1225 = i == 10'h148 ? _GEN_1224 : _GEN_1223; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1226 = ~io_inputBit ? 1'h0 : _GEN_1225; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1227 = i == 10'h265 ? _GEN_1226 : _GEN_1225; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1228 = io_inputBit | _GEN_1227; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1229 = i == 10'h265 ? _GEN_1228 : _GEN_1227; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1230 = ~io_inputBit | _GEN_1229; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1231 = i == 10'h269 ? _GEN_1230 : _GEN_1229; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1232 = io_inputBit ? 1'h0 : _GEN_1231; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1233 = i == 10'h269 ? _GEN_1232 : _GEN_1231; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1234 = ~io_inputBit ? 1'h0 : _GEN_1233; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1235 = i == 10'h26d ? _GEN_1234 : _GEN_1233; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1236 = io_inputBit | _GEN_1235; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1237 = i == 10'h26d ? _GEN_1236 : _GEN_1235; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1238 = ~io_inputBit | _GEN_1237; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1239 = i == 10'h271 ? _GEN_1238 : _GEN_1237; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1240 = io_inputBit ? 1'h0 : _GEN_1239; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1241 = i == 10'h271 ? _GEN_1240 : _GEN_1239; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1242 = ~io_inputBit ? 1'h0 : _GEN_1241; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1243 = i == 10'h275 ? _GEN_1242 : _GEN_1241; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1244 = io_inputBit | _GEN_1243; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1245 = i == 10'h275 ? _GEN_1244 : _GEN_1243; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1246 = ~io_inputBit | _GEN_1245; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1247 = i == 10'h279 ? _GEN_1246 : _GEN_1245; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1248 = io_inputBit ? 1'h0 : _GEN_1247; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1249 = i == 10'h279 ? _GEN_1248 : _GEN_1247; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1250 = ~io_inputBit ? 1'h0 : _GEN_1249; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1251 = i == 10'h27d ? _GEN_1250 : _GEN_1249; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1252 = io_inputBit | _GEN_1251; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1253 = i == 10'h27d ? _GEN_1252 : _GEN_1251; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1254 = ~io_inputBit | _GEN_1253; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1255 = i == 10'h281 ? _GEN_1254 : _GEN_1253; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1256 = io_inputBit ? 1'h0 : _GEN_1255; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1257 = i == 10'h281 ? _GEN_1256 : _GEN_1255; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1258 = ~io_inputBit ? 1'h0 : _GEN_1257; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1259 = i == 10'h285 ? _GEN_1258 : _GEN_1257; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1260 = io_inputBit | _GEN_1259; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1261 = i == 10'h285 ? _GEN_1260 : _GEN_1259; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1262 = ~io_inputBit | _GEN_1261; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1263 = i == 10'h289 ? _GEN_1262 : _GEN_1261; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1264 = io_inputBit ? 1'h0 : _GEN_1263; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1265 = i == 10'h289 ? _GEN_1264 : _GEN_1263; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1266 = ~io_inputBit ? 1'h0 : _GEN_1265; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1267 = i == 10'h28d ? _GEN_1266 : _GEN_1265; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1268 = io_inputBit | _GEN_1267; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1269 = i == 10'h28d ? _GEN_1268 : _GEN_1267; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1270 = ~io_inputBit | _GEN_1269; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1271 = i == 10'h291 ? _GEN_1270 : _GEN_1269; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1274 = io_inputBit ? 1'h0 : _GEN_415; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1275 = i == 10'h0 ? _GEN_1274 : _GEN_415; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1276 = io_inputBit ? 1'h0 : _GEN_1275; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1277 = i == 10'h4 ? _GEN_1276 : _GEN_1275; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1278 = io_inputBit ? 1'h0 : _GEN_1277; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1279 = i == 10'h9 ? _GEN_1278 : _GEN_1277; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1280 = ~io_inputBit ? 1'h0 : _GEN_1279; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1281 = i == 10'hf ? _GEN_1280 : _GEN_1279; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1282 = io_inputBit | _GEN_1281; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1283 = i == 10'h11 ? _GEN_1282 : _GEN_1281; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1284 = ~io_inputBit ? 1'h0 : _GEN_1283; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1285 = i == 10'h20 ? _GEN_1284 : _GEN_1283; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1286 = io_inputBit ? 1'h0 : _GEN_1285; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1287 = i == 10'h28 ? _GEN_1286 : _GEN_1285; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1288 = io_inputBit | _GEN_1287; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1289 = i == 10'h48 ? _GEN_1288 : _GEN_1287; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1290 = ~io_inputBit | _GEN_1289; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1291 = i == 10'h4b ? _GEN_1290 : _GEN_1289; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1292 = ~io_inputBit ? 1'h0 : _GEN_1291; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1293 = i == 10'h85 ? _GEN_1292 : _GEN_1291; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1294 = io_inputBit ? 1'h0 : _GEN_1293; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1295 = i == 10'ha4 ? _GEN_1294 : _GEN_1293; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1296 = ~io_inputBit ? 1'h0 : _GEN_1295; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1297 = i == 10'h10c ? _GEN_1296 : _GEN_1295; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1298 = io_inputBit | _GEN_1297; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1299 = i == 10'h10c ? _GEN_1298 : _GEN_1297; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1300 = ~io_inputBit | _GEN_1299; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1301 = i == 10'h10d ? _GEN_1300 : _GEN_1299; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1302 = io_inputBit ? 1'h0 : _GEN_1301; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1303 = i == 10'h10d ? _GEN_1302 : _GEN_1301; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1304 = ~io_inputBit ? 1'h0 : _GEN_1303; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1305 = i == 10'h10e ? _GEN_1304 : _GEN_1303; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1306 = io_inputBit | _GEN_1305; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1307 = i == 10'h10e ? _GEN_1306 : _GEN_1305; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1308 = ~io_inputBit | _GEN_1307; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1309 = i == 10'h10f ? _GEN_1308 : _GEN_1307; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1310 = io_inputBit ? 1'h0 : _GEN_1309; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1311 = i == 10'h10f ? _GEN_1310 : _GEN_1309; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1312 = ~io_inputBit ? 1'h0 : _GEN_1311; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1313 = i == 10'h110 ? _GEN_1312 : _GEN_1311; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1314 = io_inputBit | _GEN_1313; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1315 = i == 10'h110 ? _GEN_1314 : _GEN_1313; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1316 = ~io_inputBit | _GEN_1315; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1317 = i == 10'h111 ? _GEN_1316 : _GEN_1315; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1318 = io_inputBit ? 1'h0 : _GEN_1317; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1319 = i == 10'h111 ? _GEN_1318 : _GEN_1317; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1320 = ~io_inputBit ? 1'h0 : _GEN_1319; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1321 = i == 10'h112 ? _GEN_1320 : _GEN_1319; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1322 = io_inputBit | _GEN_1321; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1323 = i == 10'h112 ? _GEN_1322 : _GEN_1321; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1324 = ~io_inputBit | _GEN_1323; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1325 = i == 10'h113 ? _GEN_1324 : _GEN_1323; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1326 = io_inputBit ? 1'h0 : _GEN_1325; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1327 = i == 10'h113 ? _GEN_1326 : _GEN_1325; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1328 = ~io_inputBit ? 1'h0 : _GEN_1327; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1329 = i == 10'h114 ? _GEN_1328 : _GEN_1327; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1330 = io_inputBit | _GEN_1329; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1331 = i == 10'h114 ? _GEN_1330 : _GEN_1329; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1332 = ~io_inputBit | _GEN_1331; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1333 = i == 10'h115 ? _GEN_1332 : _GEN_1331; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1334 = io_inputBit ? 1'h0 : _GEN_1333; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1335 = i == 10'h115 ? _GEN_1334 : _GEN_1333; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1336 = ~io_inputBit ? 1'h0 : _GEN_1335; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1337 = i == 10'h116 ? _GEN_1336 : _GEN_1335; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1338 = io_inputBit | _GEN_1337; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1339 = i == 10'h116 ? _GEN_1338 : _GEN_1337; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1340 = ~io_inputBit | _GEN_1339; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1341 = i == 10'h117 ? _GEN_1340 : _GEN_1339; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1342 = io_inputBit ? 1'h0 : _GEN_1341; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1343 = i == 10'h117 ? _GEN_1342 : _GEN_1341; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1344 = ~io_inputBit ? 1'h0 : _GEN_1343; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1345 = i == 10'h118 ? _GEN_1344 : _GEN_1343; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1346 = io_inputBit | _GEN_1345; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1347 = i == 10'h118 ? _GEN_1346 : _GEN_1345; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1348 = ~io_inputBit | _GEN_1347; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1349 = i == 10'h119 ? _GEN_1348 : _GEN_1347; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1350 = io_inputBit ? 1'h0 : _GEN_1349; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1351 = i == 10'h119 ? _GEN_1350 : _GEN_1349; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1352 = ~io_inputBit ? 1'h0 : _GEN_1351; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1353 = i == 10'h11a ? _GEN_1352 : _GEN_1351; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1354 = io_inputBit | _GEN_1353; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1355 = i == 10'h11a ? _GEN_1354 : _GEN_1353; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1356 = ~io_inputBit | _GEN_1355; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1357 = i == 10'h11b ? _GEN_1356 : _GEN_1355; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1358 = io_inputBit ? 1'h0 : _GEN_1357; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1359 = i == 10'h11b ? _GEN_1358 : _GEN_1357; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1360 = ~io_inputBit ? 1'h0 : _GEN_1359; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1361 = i == 10'h11c ? _GEN_1360 : _GEN_1359; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1362 = io_inputBit | _GEN_1361; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1363 = i == 10'h11c ? _GEN_1362 : _GEN_1361; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1364 = ~io_inputBit | _GEN_1363; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1365 = i == 10'h11d ? _GEN_1364 : _GEN_1363; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1366 = io_inputBit ? 1'h0 : _GEN_1365; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1367 = i == 10'h11d ? _GEN_1366 : _GEN_1365; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1368 = ~io_inputBit ? 1'h0 : _GEN_1367; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1369 = i == 10'h11e ? _GEN_1368 : _GEN_1367; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1370 = io_inputBit | _GEN_1369; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1371 = i == 10'h11e ? _GEN_1370 : _GEN_1369; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1372 = ~io_inputBit | _GEN_1371; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1373 = i == 10'h11f ? _GEN_1372 : _GEN_1371; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1374 = io_inputBit ? 1'h0 : _GEN_1373; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1375 = i == 10'h11f ? _GEN_1374 : _GEN_1373; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1376 = ~io_inputBit ? 1'h0 : _GEN_1375; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1377 = i == 10'h120 ? _GEN_1376 : _GEN_1375; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1378 = io_inputBit | _GEN_1377; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1379 = i == 10'h120 ? _GEN_1378 : _GEN_1377; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1380 = ~io_inputBit | _GEN_1379; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1381 = i == 10'h121 ? _GEN_1380 : _GEN_1379; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1382 = io_inputBit ? 1'h0 : _GEN_1381; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1383 = i == 10'h121 ? _GEN_1382 : _GEN_1381; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1384 = ~io_inputBit ? 1'h0 : _GEN_1383; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1385 = i == 10'h122 ? _GEN_1384 : _GEN_1383; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1386 = io_inputBit | _GEN_1385; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1387 = i == 10'h122 ? _GEN_1386 : _GEN_1385; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1388 = ~io_inputBit | _GEN_1387; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1389 = i == 10'h123 ? _GEN_1388 : _GEN_1387; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1390 = io_inputBit ? 1'h0 : _GEN_1389; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1391 = i == 10'h123 ? _GEN_1390 : _GEN_1389; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1392 = ~io_inputBit ? 1'h0 : _GEN_1391; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1393 = i == 10'h124 ? _GEN_1392 : _GEN_1391; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1394 = io_inputBit | _GEN_1393; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1395 = i == 10'h124 ? _GEN_1394 : _GEN_1393; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1396 = io_inputBit ? 1'h0 : _GEN_1395; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1397 = i == 10'h131 ? _GEN_1396 : _GEN_1395; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1398 = io_inputBit | _GEN_1397; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1399 = i == 10'h132 ? _GEN_1398 : _GEN_1397; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1400 = io_inputBit ? 1'h0 : _GEN_1399; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1401 = i == 10'h133 ? _GEN_1400 : _GEN_1399; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1402 = io_inputBit | _GEN_1401; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1403 = i == 10'h134 ? _GEN_1402 : _GEN_1401; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1404 = io_inputBit ? 1'h0 : _GEN_1403; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1405 = i == 10'h135 ? _GEN_1404 : _GEN_1403; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1406 = io_inputBit | _GEN_1405; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1407 = i == 10'h136 ? _GEN_1406 : _GEN_1405; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1408 = io_inputBit ? 1'h0 : _GEN_1407; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1409 = i == 10'h137 ? _GEN_1408 : _GEN_1407; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1410 = io_inputBit | _GEN_1409; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1411 = i == 10'h138 ? _GEN_1410 : _GEN_1409; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1412 = io_inputBit ? 1'h0 : _GEN_1411; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1413 = i == 10'h139 ? _GEN_1412 : _GEN_1411; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1414 = io_inputBit | _GEN_1413; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1415 = i == 10'h13a ? _GEN_1414 : _GEN_1413; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1416 = io_inputBit ? 1'h0 : _GEN_1415; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1417 = i == 10'h13b ? _GEN_1416 : _GEN_1415; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1418 = io_inputBit | _GEN_1417; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1419 = i == 10'h13c ? _GEN_1418 : _GEN_1417; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1420 = io_inputBit ? 1'h0 : _GEN_1419; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1421 = i == 10'h13d ? _GEN_1420 : _GEN_1419; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1422 = io_inputBit | _GEN_1421; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1423 = i == 10'h13e ? _GEN_1422 : _GEN_1421; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1424 = io_inputBit ? 1'h0 : _GEN_1423; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1425 = i == 10'h13f ? _GEN_1424 : _GEN_1423; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1426 = io_inputBit | _GEN_1425; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1427 = i == 10'h140 ? _GEN_1426 : _GEN_1425; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1428 = io_inputBit ? 1'h0 : _GEN_1427; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1429 = i == 10'h141 ? _GEN_1428 : _GEN_1427; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1430 = io_inputBit | _GEN_1429; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1431 = i == 10'h142 ? _GEN_1430 : _GEN_1429; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1432 = io_inputBit ? 1'h0 : _GEN_1431; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1433 = i == 10'h143 ? _GEN_1432 : _GEN_1431; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1434 = io_inputBit | _GEN_1433; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1435 = i == 10'h144 ? _GEN_1434 : _GEN_1433; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1436 = io_inputBit ? 1'h0 : _GEN_1435; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1437 = i == 10'h145 ? _GEN_1436 : _GEN_1435; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1438 = io_inputBit | _GEN_1437; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1439 = i == 10'h146 ? _GEN_1438 : _GEN_1437; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1440 = io_inputBit ? 1'h0 : _GEN_1439; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1441 = i == 10'h147 ? _GEN_1440 : _GEN_1439; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1442 = io_inputBit | _GEN_1441; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1443 = i == 10'h148 ? _GEN_1442 : _GEN_1441; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1444 = io_inputBit ? 1'h0 : _GEN_1443; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1445 = i == 10'h149 ? _GEN_1444 : _GEN_1443; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1446 = ~io_inputBit | _GEN_1445; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1447 = i == 10'h263 ? _GEN_1446 : _GEN_1445; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1448 = io_inputBit ? 1'h0 : _GEN_1447; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1449 = i == 10'h263 ? _GEN_1448 : _GEN_1447; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1450 = ~io_inputBit ? 1'h0 : _GEN_1449; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1451 = i == 10'h265 ? _GEN_1450 : _GEN_1449; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1452 = io_inputBit | _GEN_1451; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1453 = i == 10'h265 ? _GEN_1452 : _GEN_1451; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1454 = ~io_inputBit | _GEN_1453; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1455 = i == 10'h267 ? _GEN_1454 : _GEN_1453; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1456 = io_inputBit ? 1'h0 : _GEN_1455; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1457 = i == 10'h267 ? _GEN_1456 : _GEN_1455; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1458 = ~io_inputBit ? 1'h0 : _GEN_1457; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1459 = i == 10'h269 ? _GEN_1458 : _GEN_1457; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1460 = io_inputBit | _GEN_1459; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1461 = i == 10'h269 ? _GEN_1460 : _GEN_1459; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1462 = ~io_inputBit | _GEN_1461; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1463 = i == 10'h26b ? _GEN_1462 : _GEN_1461; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1464 = io_inputBit ? 1'h0 : _GEN_1463; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1465 = i == 10'h26b ? _GEN_1464 : _GEN_1463; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1466 = ~io_inputBit ? 1'h0 : _GEN_1465; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1467 = i == 10'h26d ? _GEN_1466 : _GEN_1465; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1468 = io_inputBit | _GEN_1467; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1469 = i == 10'h26d ? _GEN_1468 : _GEN_1467; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1470 = ~io_inputBit | _GEN_1469; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1471 = i == 10'h26f ? _GEN_1470 : _GEN_1469; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1472 = io_inputBit ? 1'h0 : _GEN_1471; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1473 = i == 10'h26f ? _GEN_1472 : _GEN_1471; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1474 = ~io_inputBit ? 1'h0 : _GEN_1473; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1475 = i == 10'h271 ? _GEN_1474 : _GEN_1473; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1476 = io_inputBit | _GEN_1475; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1477 = i == 10'h271 ? _GEN_1476 : _GEN_1475; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1478 = ~io_inputBit | _GEN_1477; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1479 = i == 10'h273 ? _GEN_1478 : _GEN_1477; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1480 = io_inputBit ? 1'h0 : _GEN_1479; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1481 = i == 10'h273 ? _GEN_1480 : _GEN_1479; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1482 = ~io_inputBit ? 1'h0 : _GEN_1481; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1483 = i == 10'h275 ? _GEN_1482 : _GEN_1481; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1484 = io_inputBit | _GEN_1483; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1485 = i == 10'h275 ? _GEN_1484 : _GEN_1483; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1486 = ~io_inputBit | _GEN_1485; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1487 = i == 10'h277 ? _GEN_1486 : _GEN_1485; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1488 = io_inputBit ? 1'h0 : _GEN_1487; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1489 = i == 10'h277 ? _GEN_1488 : _GEN_1487; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1490 = ~io_inputBit ? 1'h0 : _GEN_1489; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1491 = i == 10'h279 ? _GEN_1490 : _GEN_1489; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1492 = io_inputBit | _GEN_1491; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1493 = i == 10'h279 ? _GEN_1492 : _GEN_1491; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1494 = ~io_inputBit | _GEN_1493; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1495 = i == 10'h27b ? _GEN_1494 : _GEN_1493; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1496 = io_inputBit ? 1'h0 : _GEN_1495; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1497 = i == 10'h27b ? _GEN_1496 : _GEN_1495; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1498 = ~io_inputBit ? 1'h0 : _GEN_1497; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1499 = i == 10'h27d ? _GEN_1498 : _GEN_1497; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1500 = io_inputBit | _GEN_1499; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1501 = i == 10'h27d ? _GEN_1500 : _GEN_1499; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1502 = ~io_inputBit | _GEN_1501; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1503 = i == 10'h27f ? _GEN_1502 : _GEN_1501; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1504 = io_inputBit ? 1'h0 : _GEN_1503; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1505 = i == 10'h27f ? _GEN_1504 : _GEN_1503; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1506 = ~io_inputBit ? 1'h0 : _GEN_1505; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1507 = i == 10'h281 ? _GEN_1506 : _GEN_1505; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1508 = io_inputBit | _GEN_1507; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1509 = i == 10'h281 ? _GEN_1508 : _GEN_1507; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1510 = ~io_inputBit | _GEN_1509; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1511 = i == 10'h283 ? _GEN_1510 : _GEN_1509; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1512 = io_inputBit ? 1'h0 : _GEN_1511; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1513 = i == 10'h283 ? _GEN_1512 : _GEN_1511; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1514 = ~io_inputBit ? 1'h0 : _GEN_1513; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1515 = i == 10'h285 ? _GEN_1514 : _GEN_1513; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1516 = io_inputBit | _GEN_1515; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1517 = i == 10'h285 ? _GEN_1516 : _GEN_1515; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1518 = ~io_inputBit | _GEN_1517; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1519 = i == 10'h287 ? _GEN_1518 : _GEN_1517; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1520 = io_inputBit ? 1'h0 : _GEN_1519; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1521 = i == 10'h287 ? _GEN_1520 : _GEN_1519; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1522 = ~io_inputBit ? 1'h0 : _GEN_1521; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1523 = i == 10'h289 ? _GEN_1522 : _GEN_1521; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1524 = io_inputBit | _GEN_1523; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1525 = i == 10'h289 ? _GEN_1524 : _GEN_1523; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1526 = ~io_inputBit | _GEN_1525; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1527 = i == 10'h28b ? _GEN_1526 : _GEN_1525; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1528 = io_inputBit ? 1'h0 : _GEN_1527; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1529 = i == 10'h28b ? _GEN_1528 : _GEN_1527; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1530 = ~io_inputBit ? 1'h0 : _GEN_1529; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1531 = i == 10'h28d ? _GEN_1530 : _GEN_1529; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1532 = io_inputBit | _GEN_1531; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1533 = i == 10'h28d ? _GEN_1532 : _GEN_1531; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1534 = ~io_inputBit | _GEN_1533; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1535 = i == 10'h28f ? _GEN_1534 : _GEN_1533; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1536 = io_inputBit ? 1'h0 : _GEN_1535; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1537 = i == 10'h28f ? _GEN_1536 : _GEN_1535; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1538 = ~io_inputBit ? 1'h0 : _GEN_1537; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1539 = i == 10'h291 ? _GEN_1538 : _GEN_1537; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1540 = io_inputBit | _GEN_1539; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1541 = i == 10'h291 ? _GEN_1540 : _GEN_1539; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1542 = ~io_inputBit | _GEN_1541; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1543 = i == 10'h293 ? _GEN_1542 : _GEN_1541; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1546 = io_inputBit ? 1'h0 : _GEN_633; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1547 = i == 10'h0 ? _GEN_1546 : _GEN_633; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1548 = io_inputBit ? 1'h0 : _GEN_1547; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1549 = i == 10'h4 ? _GEN_1548 : _GEN_1547; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1550 = io_inputBit ? 1'h0 : _GEN_1549; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1551 = i == 10'h9 ? _GEN_1550 : _GEN_1549; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1552 = ~io_inputBit ? 1'h0 : _GEN_1551; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1553 = i == 10'hf ? _GEN_1552 : _GEN_1551; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1554 = io_inputBit ? 1'h0 : _GEN_1553; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1555 = i == 10'h11 ? _GEN_1554 : _GEN_1553; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1556 = ~io_inputBit ? 1'h0 : _GEN_1555; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1557 = i == 10'h20 ? _GEN_1556 : _GEN_1555; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1558 = io_inputBit ? 1'h0 : _GEN_1557; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1559 = i == 10'h28 ? _GEN_1558 : _GEN_1557; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1560 = io_inputBit ? 1'h0 : _GEN_1559; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1561 = i == 10'h48 ? _GEN_1560 : _GEN_1559; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1562 = ~io_inputBit ? 1'h0 : _GEN_1561; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1563 = i == 10'h4b ? _GEN_1562 : _GEN_1561; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1564 = ~io_inputBit ? 1'h0 : _GEN_1563; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1565 = i == 10'h85 ? _GEN_1564 : _GEN_1563; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1566 = io_inputBit ? 1'h0 : _GEN_1565; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1567 = i == 10'ha4 ? _GEN_1566 : _GEN_1565; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1568 = ~io_inputBit | _GEN_1567; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1569 = i == 10'h10c ? _GEN_1568 : _GEN_1567; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1570 = io_inputBit ? 1'h0 : _GEN_1569; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1571 = i == 10'h10c ? _GEN_1570 : _GEN_1569; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1572 = ~io_inputBit | _GEN_1571; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1573 = i == 10'h10d ? _GEN_1572 : _GEN_1571; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1574 = io_inputBit ? 1'h0 : _GEN_1573; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1575 = i == 10'h10d ? _GEN_1574 : _GEN_1573; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1576 = ~io_inputBit | _GEN_1575; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1577 = i == 10'h10e ? _GEN_1576 : _GEN_1575; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1578 = io_inputBit ? 1'h0 : _GEN_1577; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1579 = i == 10'h10e ? _GEN_1578 : _GEN_1577; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1580 = ~io_inputBit | _GEN_1579; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1581 = i == 10'h10f ? _GEN_1580 : _GEN_1579; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1582 = io_inputBit ? 1'h0 : _GEN_1581; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1583 = i == 10'h10f ? _GEN_1582 : _GEN_1581; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1584 = ~io_inputBit | _GEN_1583; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1585 = i == 10'h110 ? _GEN_1584 : _GEN_1583; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1586 = io_inputBit ? 1'h0 : _GEN_1585; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1587 = i == 10'h110 ? _GEN_1586 : _GEN_1585; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1588 = ~io_inputBit | _GEN_1587; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1589 = i == 10'h111 ? _GEN_1588 : _GEN_1587; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1590 = io_inputBit ? 1'h0 : _GEN_1589; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1591 = i == 10'h111 ? _GEN_1590 : _GEN_1589; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1592 = ~io_inputBit | _GEN_1591; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1593 = i == 10'h112 ? _GEN_1592 : _GEN_1591; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1594 = io_inputBit ? 1'h0 : _GEN_1593; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1595 = i == 10'h112 ? _GEN_1594 : _GEN_1593; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1596 = ~io_inputBit | _GEN_1595; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1597 = i == 10'h113 ? _GEN_1596 : _GEN_1595; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1598 = io_inputBit ? 1'h0 : _GEN_1597; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1599 = i == 10'h113 ? _GEN_1598 : _GEN_1597; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1600 = ~io_inputBit | _GEN_1599; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1601 = i == 10'h114 ? _GEN_1600 : _GEN_1599; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1602 = io_inputBit ? 1'h0 : _GEN_1601; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1603 = i == 10'h114 ? _GEN_1602 : _GEN_1601; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1604 = ~io_inputBit | _GEN_1603; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1605 = i == 10'h115 ? _GEN_1604 : _GEN_1603; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1606 = io_inputBit ? 1'h0 : _GEN_1605; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1607 = i == 10'h115 ? _GEN_1606 : _GEN_1605; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1608 = ~io_inputBit | _GEN_1607; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1609 = i == 10'h116 ? _GEN_1608 : _GEN_1607; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1610 = io_inputBit ? 1'h0 : _GEN_1609; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1611 = i == 10'h116 ? _GEN_1610 : _GEN_1609; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1612 = ~io_inputBit | _GEN_1611; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1613 = i == 10'h117 ? _GEN_1612 : _GEN_1611; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1614 = io_inputBit ? 1'h0 : _GEN_1613; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1615 = i == 10'h117 ? _GEN_1614 : _GEN_1613; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1616 = ~io_inputBit | _GEN_1615; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1617 = i == 10'h118 ? _GEN_1616 : _GEN_1615; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1618 = io_inputBit ? 1'h0 : _GEN_1617; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1619 = i == 10'h118 ? _GEN_1618 : _GEN_1617; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1620 = ~io_inputBit | _GEN_1619; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1621 = i == 10'h119 ? _GEN_1620 : _GEN_1619; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1622 = io_inputBit ? 1'h0 : _GEN_1621; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1623 = i == 10'h119 ? _GEN_1622 : _GEN_1621; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1624 = ~io_inputBit | _GEN_1623; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1625 = i == 10'h11a ? _GEN_1624 : _GEN_1623; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1626 = io_inputBit ? 1'h0 : _GEN_1625; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1627 = i == 10'h11a ? _GEN_1626 : _GEN_1625; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1628 = ~io_inputBit | _GEN_1627; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1629 = i == 10'h11b ? _GEN_1628 : _GEN_1627; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1630 = io_inputBit ? 1'h0 : _GEN_1629; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1631 = i == 10'h11b ? _GEN_1630 : _GEN_1629; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1632 = ~io_inputBit | _GEN_1631; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1633 = i == 10'h11c ? _GEN_1632 : _GEN_1631; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1634 = io_inputBit ? 1'h0 : _GEN_1633; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1635 = i == 10'h11c ? _GEN_1634 : _GEN_1633; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1636 = ~io_inputBit | _GEN_1635; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1637 = i == 10'h11d ? _GEN_1636 : _GEN_1635; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1638 = io_inputBit ? 1'h0 : _GEN_1637; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1639 = i == 10'h11d ? _GEN_1638 : _GEN_1637; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1640 = ~io_inputBit | _GEN_1639; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1641 = i == 10'h11e ? _GEN_1640 : _GEN_1639; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1642 = io_inputBit ? 1'h0 : _GEN_1641; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1643 = i == 10'h11e ? _GEN_1642 : _GEN_1641; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1644 = ~io_inputBit | _GEN_1643; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1645 = i == 10'h11f ? _GEN_1644 : _GEN_1643; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1646 = io_inputBit ? 1'h0 : _GEN_1645; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1647 = i == 10'h11f ? _GEN_1646 : _GEN_1645; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1648 = ~io_inputBit | _GEN_1647; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1649 = i == 10'h120 ? _GEN_1648 : _GEN_1647; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1650 = io_inputBit ? 1'h0 : _GEN_1649; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1651 = i == 10'h120 ? _GEN_1650 : _GEN_1649; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1652 = ~io_inputBit | _GEN_1651; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1653 = i == 10'h121 ? _GEN_1652 : _GEN_1651; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1654 = io_inputBit ? 1'h0 : _GEN_1653; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1655 = i == 10'h121 ? _GEN_1654 : _GEN_1653; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1656 = ~io_inputBit | _GEN_1655; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1657 = i == 10'h122 ? _GEN_1656 : _GEN_1655; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1658 = io_inputBit ? 1'h0 : _GEN_1657; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1659 = i == 10'h122 ? _GEN_1658 : _GEN_1657; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1660 = ~io_inputBit | _GEN_1659; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1661 = i == 10'h123 ? _GEN_1660 : _GEN_1659; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1662 = io_inputBit ? 1'h0 : _GEN_1661; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1663 = i == 10'h123 ? _GEN_1662 : _GEN_1661; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1664 = ~io_inputBit | _GEN_1663; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1665 = i == 10'h124 ? _GEN_1664 : _GEN_1663; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1666 = io_inputBit ? 1'h0 : _GEN_1665; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1667 = i == 10'h124 ? _GEN_1666 : _GEN_1665; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1668 = ~io_inputBit ? 1'h0 : _GEN_1667; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1669 = i == 10'h263 ? _GEN_1668 : _GEN_1667; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1670 = io_inputBit | _GEN_1669; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1671 = i == 10'h263 ? _GEN_1670 : _GEN_1669; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1672 = ~io_inputBit | _GEN_1671; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1673 = i == 10'h264 ? _GEN_1672 : _GEN_1671; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1674 = io_inputBit ? 1'h0 : _GEN_1673; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1675 = i == 10'h264 ? _GEN_1674 : _GEN_1673; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1676 = ~io_inputBit ? 1'h0 : _GEN_1675; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1677 = i == 10'h265 ? _GEN_1676 : _GEN_1675; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1678 = io_inputBit | _GEN_1677; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1679 = i == 10'h265 ? _GEN_1678 : _GEN_1677; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1680 = ~io_inputBit | _GEN_1679; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1681 = i == 10'h266 ? _GEN_1680 : _GEN_1679; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1682 = io_inputBit ? 1'h0 : _GEN_1681; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1683 = i == 10'h266 ? _GEN_1682 : _GEN_1681; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1684 = ~io_inputBit ? 1'h0 : _GEN_1683; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1685 = i == 10'h267 ? _GEN_1684 : _GEN_1683; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1686 = io_inputBit | _GEN_1685; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1687 = i == 10'h267 ? _GEN_1686 : _GEN_1685; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1688 = ~io_inputBit | _GEN_1687; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1689 = i == 10'h268 ? _GEN_1688 : _GEN_1687; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1690 = io_inputBit ? 1'h0 : _GEN_1689; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1691 = i == 10'h268 ? _GEN_1690 : _GEN_1689; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1692 = ~io_inputBit ? 1'h0 : _GEN_1691; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1693 = i == 10'h269 ? _GEN_1692 : _GEN_1691; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1694 = io_inputBit | _GEN_1693; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1695 = i == 10'h269 ? _GEN_1694 : _GEN_1693; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1696 = ~io_inputBit | _GEN_1695; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1697 = i == 10'h26a ? _GEN_1696 : _GEN_1695; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1698 = io_inputBit ? 1'h0 : _GEN_1697; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1699 = i == 10'h26a ? _GEN_1698 : _GEN_1697; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1700 = ~io_inputBit ? 1'h0 : _GEN_1699; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1701 = i == 10'h26b ? _GEN_1700 : _GEN_1699; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1702 = io_inputBit | _GEN_1701; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1703 = i == 10'h26b ? _GEN_1702 : _GEN_1701; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1704 = ~io_inputBit | _GEN_1703; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1705 = i == 10'h26c ? _GEN_1704 : _GEN_1703; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1706 = io_inputBit ? 1'h0 : _GEN_1705; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1707 = i == 10'h26c ? _GEN_1706 : _GEN_1705; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1708 = ~io_inputBit ? 1'h0 : _GEN_1707; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1709 = i == 10'h26d ? _GEN_1708 : _GEN_1707; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1710 = io_inputBit | _GEN_1709; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1711 = i == 10'h26d ? _GEN_1710 : _GEN_1709; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1712 = ~io_inputBit | _GEN_1711; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1713 = i == 10'h26e ? _GEN_1712 : _GEN_1711; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1714 = io_inputBit ? 1'h0 : _GEN_1713; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1715 = i == 10'h26e ? _GEN_1714 : _GEN_1713; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1716 = ~io_inputBit ? 1'h0 : _GEN_1715; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1717 = i == 10'h26f ? _GEN_1716 : _GEN_1715; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1718 = io_inputBit | _GEN_1717; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1719 = i == 10'h26f ? _GEN_1718 : _GEN_1717; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1720 = ~io_inputBit | _GEN_1719; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1721 = i == 10'h270 ? _GEN_1720 : _GEN_1719; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1722 = io_inputBit ? 1'h0 : _GEN_1721; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1723 = i == 10'h270 ? _GEN_1722 : _GEN_1721; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1724 = ~io_inputBit ? 1'h0 : _GEN_1723; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1725 = i == 10'h271 ? _GEN_1724 : _GEN_1723; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1726 = io_inputBit | _GEN_1725; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1727 = i == 10'h271 ? _GEN_1726 : _GEN_1725; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1728 = ~io_inputBit | _GEN_1727; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1729 = i == 10'h272 ? _GEN_1728 : _GEN_1727; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1730 = io_inputBit ? 1'h0 : _GEN_1729; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1731 = i == 10'h272 ? _GEN_1730 : _GEN_1729; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1732 = ~io_inputBit ? 1'h0 : _GEN_1731; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1733 = i == 10'h273 ? _GEN_1732 : _GEN_1731; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1734 = io_inputBit | _GEN_1733; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1735 = i == 10'h273 ? _GEN_1734 : _GEN_1733; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1736 = ~io_inputBit | _GEN_1735; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1737 = i == 10'h274 ? _GEN_1736 : _GEN_1735; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1738 = io_inputBit ? 1'h0 : _GEN_1737; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1739 = i == 10'h274 ? _GEN_1738 : _GEN_1737; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1740 = ~io_inputBit ? 1'h0 : _GEN_1739; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1741 = i == 10'h275 ? _GEN_1740 : _GEN_1739; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1742 = io_inputBit | _GEN_1741; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1743 = i == 10'h275 ? _GEN_1742 : _GEN_1741; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1744 = ~io_inputBit | _GEN_1743; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1745 = i == 10'h276 ? _GEN_1744 : _GEN_1743; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1746 = io_inputBit ? 1'h0 : _GEN_1745; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1747 = i == 10'h276 ? _GEN_1746 : _GEN_1745; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1748 = ~io_inputBit ? 1'h0 : _GEN_1747; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1749 = i == 10'h277 ? _GEN_1748 : _GEN_1747; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1750 = io_inputBit | _GEN_1749; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1751 = i == 10'h277 ? _GEN_1750 : _GEN_1749; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1752 = ~io_inputBit | _GEN_1751; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1753 = i == 10'h278 ? _GEN_1752 : _GEN_1751; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1754 = io_inputBit ? 1'h0 : _GEN_1753; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1755 = i == 10'h278 ? _GEN_1754 : _GEN_1753; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1756 = ~io_inputBit ? 1'h0 : _GEN_1755; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1757 = i == 10'h279 ? _GEN_1756 : _GEN_1755; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1758 = io_inputBit | _GEN_1757; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1759 = i == 10'h279 ? _GEN_1758 : _GEN_1757; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1760 = ~io_inputBit | _GEN_1759; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1761 = i == 10'h27a ? _GEN_1760 : _GEN_1759; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1762 = io_inputBit ? 1'h0 : _GEN_1761; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1763 = i == 10'h27a ? _GEN_1762 : _GEN_1761; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1764 = ~io_inputBit ? 1'h0 : _GEN_1763; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1765 = i == 10'h27b ? _GEN_1764 : _GEN_1763; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1766 = io_inputBit | _GEN_1765; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1767 = i == 10'h27b ? _GEN_1766 : _GEN_1765; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1768 = ~io_inputBit | _GEN_1767; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1769 = i == 10'h27c ? _GEN_1768 : _GEN_1767; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1770 = io_inputBit ? 1'h0 : _GEN_1769; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1771 = i == 10'h27c ? _GEN_1770 : _GEN_1769; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1772 = ~io_inputBit ? 1'h0 : _GEN_1771; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1773 = i == 10'h27d ? _GEN_1772 : _GEN_1771; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1774 = io_inputBit | _GEN_1773; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1775 = i == 10'h27d ? _GEN_1774 : _GEN_1773; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1776 = ~io_inputBit | _GEN_1775; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1777 = i == 10'h27e ? _GEN_1776 : _GEN_1775; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1778 = io_inputBit ? 1'h0 : _GEN_1777; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1779 = i == 10'h27e ? _GEN_1778 : _GEN_1777; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1780 = ~io_inputBit ? 1'h0 : _GEN_1779; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1781 = i == 10'h27f ? _GEN_1780 : _GEN_1779; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1782 = io_inputBit | _GEN_1781; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1783 = i == 10'h27f ? _GEN_1782 : _GEN_1781; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1784 = ~io_inputBit | _GEN_1783; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1785 = i == 10'h280 ? _GEN_1784 : _GEN_1783; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1786 = io_inputBit ? 1'h0 : _GEN_1785; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1787 = i == 10'h280 ? _GEN_1786 : _GEN_1785; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1788 = ~io_inputBit ? 1'h0 : _GEN_1787; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1789 = i == 10'h281 ? _GEN_1788 : _GEN_1787; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1790 = io_inputBit | _GEN_1789; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1791 = i == 10'h281 ? _GEN_1790 : _GEN_1789; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1792 = ~io_inputBit | _GEN_1791; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1793 = i == 10'h282 ? _GEN_1792 : _GEN_1791; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1794 = io_inputBit ? 1'h0 : _GEN_1793; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1795 = i == 10'h282 ? _GEN_1794 : _GEN_1793; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1796 = ~io_inputBit ? 1'h0 : _GEN_1795; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1797 = i == 10'h283 ? _GEN_1796 : _GEN_1795; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1798 = io_inputBit | _GEN_1797; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1799 = i == 10'h283 ? _GEN_1798 : _GEN_1797; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1800 = ~io_inputBit | _GEN_1799; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1801 = i == 10'h284 ? _GEN_1800 : _GEN_1799; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1802 = io_inputBit ? 1'h0 : _GEN_1801; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1803 = i == 10'h284 ? _GEN_1802 : _GEN_1801; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1804 = ~io_inputBit ? 1'h0 : _GEN_1803; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1805 = i == 10'h285 ? _GEN_1804 : _GEN_1803; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1806 = io_inputBit | _GEN_1805; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1807 = i == 10'h285 ? _GEN_1806 : _GEN_1805; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1808 = ~io_inputBit | _GEN_1807; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1809 = i == 10'h286 ? _GEN_1808 : _GEN_1807; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1810 = io_inputBit ? 1'h0 : _GEN_1809; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1811 = i == 10'h286 ? _GEN_1810 : _GEN_1809; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1812 = ~io_inputBit ? 1'h0 : _GEN_1811; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1813 = i == 10'h287 ? _GEN_1812 : _GEN_1811; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1814 = io_inputBit | _GEN_1813; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1815 = i == 10'h287 ? _GEN_1814 : _GEN_1813; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1816 = ~io_inputBit | _GEN_1815; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1817 = i == 10'h288 ? _GEN_1816 : _GEN_1815; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1818 = io_inputBit ? 1'h0 : _GEN_1817; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1819 = i == 10'h288 ? _GEN_1818 : _GEN_1817; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1820 = ~io_inputBit ? 1'h0 : _GEN_1819; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1821 = i == 10'h289 ? _GEN_1820 : _GEN_1819; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1822 = io_inputBit | _GEN_1821; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1823 = i == 10'h289 ? _GEN_1822 : _GEN_1821; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1824 = ~io_inputBit | _GEN_1823; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1825 = i == 10'h28a ? _GEN_1824 : _GEN_1823; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1826 = io_inputBit ? 1'h0 : _GEN_1825; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1827 = i == 10'h28a ? _GEN_1826 : _GEN_1825; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1828 = ~io_inputBit ? 1'h0 : _GEN_1827; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1829 = i == 10'h28b ? _GEN_1828 : _GEN_1827; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1830 = io_inputBit | _GEN_1829; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1831 = i == 10'h28b ? _GEN_1830 : _GEN_1829; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1832 = ~io_inputBit | _GEN_1831; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1833 = i == 10'h28c ? _GEN_1832 : _GEN_1831; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1834 = io_inputBit ? 1'h0 : _GEN_1833; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1835 = i == 10'h28c ? _GEN_1834 : _GEN_1833; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1836 = ~io_inputBit ? 1'h0 : _GEN_1835; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1837 = i == 10'h28d ? _GEN_1836 : _GEN_1835; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1838 = io_inputBit | _GEN_1837; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1839 = i == 10'h28d ? _GEN_1838 : _GEN_1837; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1840 = ~io_inputBit | _GEN_1839; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1841 = i == 10'h28e ? _GEN_1840 : _GEN_1839; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1842 = io_inputBit ? 1'h0 : _GEN_1841; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1843 = i == 10'h28e ? _GEN_1842 : _GEN_1841; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1844 = ~io_inputBit ? 1'h0 : _GEN_1843; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1845 = i == 10'h28f ? _GEN_1844 : _GEN_1843; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1846 = io_inputBit | _GEN_1845; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1847 = i == 10'h28f ? _GEN_1846 : _GEN_1845; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1848 = ~io_inputBit | _GEN_1847; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1849 = i == 10'h290 ? _GEN_1848 : _GEN_1847; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1850 = io_inputBit ? 1'h0 : _GEN_1849; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1851 = i == 10'h290 ? _GEN_1850 : _GEN_1849; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1852 = ~io_inputBit ? 1'h0 : _GEN_1851; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1853 = i == 10'h291 ? _GEN_1852 : _GEN_1851; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1854 = io_inputBit | _GEN_1853; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1855 = i == 10'h291 ? _GEN_1854 : _GEN_1853; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1856 = ~io_inputBit | _GEN_1855; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1857 = i == 10'h292 ? _GEN_1856 : _GEN_1855; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1858 = io_inputBit ? 1'h0 : _GEN_1857; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1859 = i == 10'h292 ? _GEN_1858 : _GEN_1857; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1860 = ~io_inputBit ? 1'h0 : _GEN_1859; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1861 = i == 10'h293 ? _GEN_1860 : _GEN_1859; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1862 = io_inputBit | _GEN_1861; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1863 = i == 10'h293 ? _GEN_1862 : _GEN_1861; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1864 = ~io_inputBit | _GEN_1863; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1865 = i == 10'h294 ? _GEN_1864 : _GEN_1863; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1868 = io_inputBit ? 1'h0 : _GEN_851; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1869 = i == 10'h0 ? _GEN_1868 : _GEN_851; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1870 = io_inputBit ? 1'h0 : _GEN_1869; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1871 = i == 10'h4 ? _GEN_1870 : _GEN_1869; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1872 = io_inputBit ? 1'h0 : _GEN_1871; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1873 = i == 10'h9 ? _GEN_1872 : _GEN_1871; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1874 = ~io_inputBit ? 1'h0 : _GEN_1873; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1875 = i == 10'hf ? _GEN_1874 : _GEN_1873; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1876 = io_inputBit ? 1'h0 : _GEN_1875; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1877 = i == 10'h11 ? _GEN_1876 : _GEN_1875; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1878 = ~io_inputBit ? 1'h0 : _GEN_1877; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1879 = i == 10'h20 ? _GEN_1878 : _GEN_1877; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1880 = io_inputBit ? 1'h0 : _GEN_1879; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1881 = i == 10'h28 ? _GEN_1880 : _GEN_1879; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1882 = io_inputBit ? 1'h0 : _GEN_1881; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1883 = i == 10'h48 ? _GEN_1882 : _GEN_1881; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1884 = ~io_inputBit ? 1'h0 : _GEN_1883; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1885 = i == 10'h4b ? _GEN_1884 : _GEN_1883; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1886 = io_inputBit ? 1'h0 : _GEN_1885; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1887 = i == 10'ha4 ? _GEN_1886 : _GEN_1885; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1888 = ~io_inputBit ? 1'h0 : _GEN_1887; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1889 = i == 10'h10b ? _GEN_1888 : _GEN_1887; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1890 = io_inputBit ? 1'h0 : _GEN_1889; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1891 = i == 10'h124 ? _GEN_1890 : _GEN_1889; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1892 = ~io_inputBit ? 1'h0 : _GEN_1891; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1893 = i == 10'h218 ? _GEN_1892 : _GEN_1891; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1894 = io_inputBit | _GEN_1893; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1895 = i == 10'h218 ? _GEN_1894 : _GEN_1893; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1896 = ~io_inputBit ? 1'h0 : _GEN_1895; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1897 = i == 10'h219 ? _GEN_1896 : _GEN_1895; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1898 = io_inputBit | _GEN_1897; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1899 = i == 10'h219 ? _GEN_1898 : _GEN_1897; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1900 = ~io_inputBit ? 1'h0 : _GEN_1899; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1901 = i == 10'h21a ? _GEN_1900 : _GEN_1899; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1902 = io_inputBit | _GEN_1901; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1903 = i == 10'h21a ? _GEN_1902 : _GEN_1901; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1904 = ~io_inputBit ? 1'h0 : _GEN_1903; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1905 = i == 10'h21b ? _GEN_1904 : _GEN_1903; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1906 = io_inputBit | _GEN_1905; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1907 = i == 10'h21b ? _GEN_1906 : _GEN_1905; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1908 = ~io_inputBit ? 1'h0 : _GEN_1907; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1909 = i == 10'h21c ? _GEN_1908 : _GEN_1907; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1910 = io_inputBit | _GEN_1909; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1911 = i == 10'h21c ? _GEN_1910 : _GEN_1909; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1912 = ~io_inputBit ? 1'h0 : _GEN_1911; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1913 = i == 10'h21d ? _GEN_1912 : _GEN_1911; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1914 = io_inputBit | _GEN_1913; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1915 = i == 10'h21d ? _GEN_1914 : _GEN_1913; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1916 = ~io_inputBit ? 1'h0 : _GEN_1915; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1917 = i == 10'h21e ? _GEN_1916 : _GEN_1915; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1918 = io_inputBit | _GEN_1917; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1919 = i == 10'h21e ? _GEN_1918 : _GEN_1917; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1920 = ~io_inputBit ? 1'h0 : _GEN_1919; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1921 = i == 10'h21f ? _GEN_1920 : _GEN_1919; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1922 = io_inputBit | _GEN_1921; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1923 = i == 10'h21f ? _GEN_1922 : _GEN_1921; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1924 = ~io_inputBit ? 1'h0 : _GEN_1923; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1925 = i == 10'h220 ? _GEN_1924 : _GEN_1923; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1926 = io_inputBit | _GEN_1925; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1927 = i == 10'h220 ? _GEN_1926 : _GEN_1925; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1928 = ~io_inputBit ? 1'h0 : _GEN_1927; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1929 = i == 10'h221 ? _GEN_1928 : _GEN_1927; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1930 = io_inputBit | _GEN_1929; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1931 = i == 10'h221 ? _GEN_1930 : _GEN_1929; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1932 = ~io_inputBit ? 1'h0 : _GEN_1931; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1933 = i == 10'h222 ? _GEN_1932 : _GEN_1931; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1934 = io_inputBit | _GEN_1933; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1935 = i == 10'h222 ? _GEN_1934 : _GEN_1933; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1936 = ~io_inputBit ? 1'h0 : _GEN_1935; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1937 = i == 10'h223 ? _GEN_1936 : _GEN_1935; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1938 = io_inputBit | _GEN_1937; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1939 = i == 10'h223 ? _GEN_1938 : _GEN_1937; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1940 = ~io_inputBit ? 1'h0 : _GEN_1939; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1941 = i == 10'h224 ? _GEN_1940 : _GEN_1939; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1942 = io_inputBit | _GEN_1941; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1943 = i == 10'h224 ? _GEN_1942 : _GEN_1941; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1944 = ~io_inputBit ? 1'h0 : _GEN_1943; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1945 = i == 10'h225 ? _GEN_1944 : _GEN_1943; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1946 = io_inputBit | _GEN_1945; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1947 = i == 10'h225 ? _GEN_1946 : _GEN_1945; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1948 = ~io_inputBit ? 1'h0 : _GEN_1947; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1949 = i == 10'h226 ? _GEN_1948 : _GEN_1947; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1950 = io_inputBit | _GEN_1949; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1951 = i == 10'h226 ? _GEN_1950 : _GEN_1949; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1952 = ~io_inputBit ? 1'h0 : _GEN_1951; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1953 = i == 10'h227 ? _GEN_1952 : _GEN_1951; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1954 = io_inputBit | _GEN_1953; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1955 = i == 10'h227 ? _GEN_1954 : _GEN_1953; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1956 = ~io_inputBit ? 1'h0 : _GEN_1955; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1957 = i == 10'h228 ? _GEN_1956 : _GEN_1955; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1958 = io_inputBit | _GEN_1957; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1959 = i == 10'h228 ? _GEN_1958 : _GEN_1957; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1960 = ~io_inputBit ? 1'h0 : _GEN_1959; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1961 = i == 10'h229 ? _GEN_1960 : _GEN_1959; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1962 = io_inputBit | _GEN_1961; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1963 = i == 10'h229 ? _GEN_1962 : _GEN_1961; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1964 = ~io_inputBit ? 1'h0 : _GEN_1963; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1965 = i == 10'h22a ? _GEN_1964 : _GEN_1963; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1966 = io_inputBit | _GEN_1965; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1967 = i == 10'h22a ? _GEN_1966 : _GEN_1965; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1968 = ~io_inputBit ? 1'h0 : _GEN_1967; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1969 = i == 10'h22b ? _GEN_1968 : _GEN_1967; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1970 = io_inputBit | _GEN_1969; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1971 = i == 10'h22b ? _GEN_1970 : _GEN_1969; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1972 = ~io_inputBit ? 1'h0 : _GEN_1971; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1973 = i == 10'h22c ? _GEN_1972 : _GEN_1971; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1974 = io_inputBit | _GEN_1973; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1975 = i == 10'h22c ? _GEN_1974 : _GEN_1973; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1976 = ~io_inputBit ? 1'h0 : _GEN_1975; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1977 = i == 10'h22d ? _GEN_1976 : _GEN_1975; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1978 = io_inputBit | _GEN_1977; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1979 = i == 10'h22d ? _GEN_1978 : _GEN_1977; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1980 = ~io_inputBit ? 1'h0 : _GEN_1979; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1981 = i == 10'h22e ? _GEN_1980 : _GEN_1979; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1982 = io_inputBit | _GEN_1981; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1983 = i == 10'h22e ? _GEN_1982 : _GEN_1981; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1984 = ~io_inputBit ? 1'h0 : _GEN_1983; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1985 = i == 10'h22f ? _GEN_1984 : _GEN_1983; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1986 = io_inputBit | _GEN_1985; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1987 = i == 10'h22f ? _GEN_1986 : _GEN_1985; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1988 = ~io_inputBit ? 1'h0 : _GEN_1987; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1989 = i == 10'h230 ? _GEN_1988 : _GEN_1987; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1990 = io_inputBit | _GEN_1989; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1991 = i == 10'h230 ? _GEN_1990 : _GEN_1989; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1992 = ~io_inputBit ? 1'h0 : _GEN_1991; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1993 = i == 10'h231 ? _GEN_1992 : _GEN_1991; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1994 = io_inputBit | _GEN_1993; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1995 = i == 10'h231 ? _GEN_1994 : _GEN_1993; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1996 = ~io_inputBit ? 1'h0 : _GEN_1995; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1997 = i == 10'h232 ? _GEN_1996 : _GEN_1995; // @[lut_mem_online.scala 247:34]
  wire  _GEN_1998 = io_inputBit | _GEN_1997; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_1999 = i == 10'h232 ? _GEN_1998 : _GEN_1997; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2000 = ~io_inputBit ? 1'h0 : _GEN_1999; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2001 = i == 10'h233 ? _GEN_2000 : _GEN_1999; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2002 = io_inputBit | _GEN_2001; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2003 = i == 10'h233 ? _GEN_2002 : _GEN_2001; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2004 = ~io_inputBit ? 1'h0 : _GEN_2003; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2005 = i == 10'h234 ? _GEN_2004 : _GEN_2003; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2006 = io_inputBit | _GEN_2005; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2007 = i == 10'h234 ? _GEN_2006 : _GEN_2005; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2008 = ~io_inputBit ? 1'h0 : _GEN_2007; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2009 = i == 10'h235 ? _GEN_2008 : _GEN_2007; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2010 = io_inputBit | _GEN_2009; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2011 = i == 10'h235 ? _GEN_2010 : _GEN_2009; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2012 = ~io_inputBit ? 1'h0 : _GEN_2011; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2013 = i == 10'h236 ? _GEN_2012 : _GEN_2011; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2014 = io_inputBit | _GEN_2013; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2015 = i == 10'h236 ? _GEN_2014 : _GEN_2013; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2016 = ~io_inputBit ? 1'h0 : _GEN_2015; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2017 = i == 10'h237 ? _GEN_2016 : _GEN_2015; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2018 = io_inputBit | _GEN_2017; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2019 = i == 10'h237 ? _GEN_2018 : _GEN_2017; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2020 = ~io_inputBit ? 1'h0 : _GEN_2019; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2021 = i == 10'h238 ? _GEN_2020 : _GEN_2019; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2022 = io_inputBit | _GEN_2021; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2023 = i == 10'h238 ? _GEN_2022 : _GEN_2021; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2024 = ~io_inputBit ? 1'h0 : _GEN_2023; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2025 = i == 10'h239 ? _GEN_2024 : _GEN_2023; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2026 = io_inputBit | _GEN_2025; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2027 = i == 10'h239 ? _GEN_2026 : _GEN_2025; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2028 = ~io_inputBit ? 1'h0 : _GEN_2027; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2029 = i == 10'h23a ? _GEN_2028 : _GEN_2027; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2030 = io_inputBit | _GEN_2029; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2031 = i == 10'h23a ? _GEN_2030 : _GEN_2029; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2032 = ~io_inputBit ? 1'h0 : _GEN_2031; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2033 = i == 10'h23b ? _GEN_2032 : _GEN_2031; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2034 = io_inputBit | _GEN_2033; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2035 = i == 10'h23b ? _GEN_2034 : _GEN_2033; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2036 = ~io_inputBit ? 1'h0 : _GEN_2035; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2037 = i == 10'h23c ? _GEN_2036 : _GEN_2035; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2038 = io_inputBit | _GEN_2037; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2039 = i == 10'h23c ? _GEN_2038 : _GEN_2037; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2040 = ~io_inputBit ? 1'h0 : _GEN_2039; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2041 = i == 10'h23d ? _GEN_2040 : _GEN_2039; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2042 = io_inputBit | _GEN_2041; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2043 = i == 10'h23d ? _GEN_2042 : _GEN_2041; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2044 = ~io_inputBit ? 1'h0 : _GEN_2043; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2045 = i == 10'h23e ? _GEN_2044 : _GEN_2043; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2046 = io_inputBit | _GEN_2045; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2047 = i == 10'h23e ? _GEN_2046 : _GEN_2045; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2048 = ~io_inputBit ? 1'h0 : _GEN_2047; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2049 = i == 10'h23f ? _GEN_2048 : _GEN_2047; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2050 = io_inputBit | _GEN_2049; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2051 = i == 10'h23f ? _GEN_2050 : _GEN_2049; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2052 = ~io_inputBit ? 1'h0 : _GEN_2051; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2053 = i == 10'h240 ? _GEN_2052 : _GEN_2051; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2054 = io_inputBit | _GEN_2053; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2055 = i == 10'h240 ? _GEN_2054 : _GEN_2053; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2056 = ~io_inputBit ? 1'h0 : _GEN_2055; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2057 = i == 10'h241 ? _GEN_2056 : _GEN_2055; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2058 = io_inputBit | _GEN_2057; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2059 = i == 10'h241 ? _GEN_2058 : _GEN_2057; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2060 = ~io_inputBit ? 1'h0 : _GEN_2059; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2061 = i == 10'h242 ? _GEN_2060 : _GEN_2059; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2062 = io_inputBit | _GEN_2061; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2063 = i == 10'h242 ? _GEN_2062 : _GEN_2061; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2064 = ~io_inputBit ? 1'h0 : _GEN_2063; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2065 = i == 10'h243 ? _GEN_2064 : _GEN_2063; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2066 = io_inputBit | _GEN_2065; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2067 = i == 10'h243 ? _GEN_2066 : _GEN_2065; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2068 = ~io_inputBit ? 1'h0 : _GEN_2067; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2069 = i == 10'h244 ? _GEN_2068 : _GEN_2067; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2070 = io_inputBit | _GEN_2069; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2071 = i == 10'h244 ? _GEN_2070 : _GEN_2069; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2072 = ~io_inputBit ? 1'h0 : _GEN_2071; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2073 = i == 10'h245 ? _GEN_2072 : _GEN_2071; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2074 = io_inputBit | _GEN_2073; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2075 = i == 10'h245 ? _GEN_2074 : _GEN_2073; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2076 = ~io_inputBit ? 1'h0 : _GEN_2075; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2077 = i == 10'h246 ? _GEN_2076 : _GEN_2075; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2078 = io_inputBit | _GEN_2077; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2079 = i == 10'h246 ? _GEN_2078 : _GEN_2077; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2080 = ~io_inputBit ? 1'h0 : _GEN_2079; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2081 = i == 10'h247 ? _GEN_2080 : _GEN_2079; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2082 = io_inputBit | _GEN_2081; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2083 = i == 10'h247 ? _GEN_2082 : _GEN_2081; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2084 = ~io_inputBit ? 1'h0 : _GEN_2083; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2085 = i == 10'h248 ? _GEN_2084 : _GEN_2083; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2086 = io_inputBit | _GEN_2085; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2087 = i == 10'h248 ? _GEN_2086 : _GEN_2085; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2088 = ~io_inputBit ? 1'h0 : _GEN_2087; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2089 = i == 10'h249 ? _GEN_2088 : _GEN_2087; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2090 = io_inputBit | _GEN_2089; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2091 = i == 10'h249 ? _GEN_2090 : _GEN_2089; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2092 = ~io_inputBit ? 1'h0 : _GEN_2091; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2093 = i == 10'h263 ? _GEN_2092 : _GEN_2091; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2094 = io_inputBit | _GEN_2093; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2095 = i == 10'h263 ? _GEN_2094 : _GEN_2093; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2096 = ~io_inputBit ? 1'h0 : _GEN_2095; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2097 = i == 10'h264 ? _GEN_2096 : _GEN_2095; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2098 = io_inputBit | _GEN_2097; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2099 = i == 10'h264 ? _GEN_2098 : _GEN_2097; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2100 = ~io_inputBit ? 1'h0 : _GEN_2099; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2101 = i == 10'h265 ? _GEN_2100 : _GEN_2099; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2102 = io_inputBit | _GEN_2101; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2103 = i == 10'h265 ? _GEN_2102 : _GEN_2101; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2104 = ~io_inputBit ? 1'h0 : _GEN_2103; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2105 = i == 10'h266 ? _GEN_2104 : _GEN_2103; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2106 = io_inputBit | _GEN_2105; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2107 = i == 10'h266 ? _GEN_2106 : _GEN_2105; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2108 = ~io_inputBit ? 1'h0 : _GEN_2107; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2109 = i == 10'h267 ? _GEN_2108 : _GEN_2107; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2110 = io_inputBit | _GEN_2109; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2111 = i == 10'h267 ? _GEN_2110 : _GEN_2109; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2112 = ~io_inputBit ? 1'h0 : _GEN_2111; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2113 = i == 10'h268 ? _GEN_2112 : _GEN_2111; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2114 = io_inputBit | _GEN_2113; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2115 = i == 10'h268 ? _GEN_2114 : _GEN_2113; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2116 = ~io_inputBit ? 1'h0 : _GEN_2115; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2117 = i == 10'h269 ? _GEN_2116 : _GEN_2115; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2118 = io_inputBit | _GEN_2117; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2119 = i == 10'h269 ? _GEN_2118 : _GEN_2117; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2120 = ~io_inputBit ? 1'h0 : _GEN_2119; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2121 = i == 10'h26a ? _GEN_2120 : _GEN_2119; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2122 = io_inputBit | _GEN_2121; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2123 = i == 10'h26a ? _GEN_2122 : _GEN_2121; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2124 = ~io_inputBit ? 1'h0 : _GEN_2123; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2125 = i == 10'h26b ? _GEN_2124 : _GEN_2123; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2126 = io_inputBit | _GEN_2125; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2127 = i == 10'h26b ? _GEN_2126 : _GEN_2125; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2128 = ~io_inputBit ? 1'h0 : _GEN_2127; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2129 = i == 10'h26c ? _GEN_2128 : _GEN_2127; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2130 = io_inputBit | _GEN_2129; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2131 = i == 10'h26c ? _GEN_2130 : _GEN_2129; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2132 = ~io_inputBit ? 1'h0 : _GEN_2131; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2133 = i == 10'h26d ? _GEN_2132 : _GEN_2131; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2134 = io_inputBit | _GEN_2133; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2135 = i == 10'h26d ? _GEN_2134 : _GEN_2133; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2136 = ~io_inputBit ? 1'h0 : _GEN_2135; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2137 = i == 10'h26e ? _GEN_2136 : _GEN_2135; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2138 = io_inputBit | _GEN_2137; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2139 = i == 10'h26e ? _GEN_2138 : _GEN_2137; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2140 = ~io_inputBit ? 1'h0 : _GEN_2139; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2141 = i == 10'h26f ? _GEN_2140 : _GEN_2139; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2142 = io_inputBit | _GEN_2141; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2143 = i == 10'h26f ? _GEN_2142 : _GEN_2141; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2144 = ~io_inputBit ? 1'h0 : _GEN_2143; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2145 = i == 10'h270 ? _GEN_2144 : _GEN_2143; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2146 = io_inputBit | _GEN_2145; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2147 = i == 10'h270 ? _GEN_2146 : _GEN_2145; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2148 = ~io_inputBit ? 1'h0 : _GEN_2147; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2149 = i == 10'h271 ? _GEN_2148 : _GEN_2147; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2150 = io_inputBit | _GEN_2149; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2151 = i == 10'h271 ? _GEN_2150 : _GEN_2149; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2152 = ~io_inputBit ? 1'h0 : _GEN_2151; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2153 = i == 10'h272 ? _GEN_2152 : _GEN_2151; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2154 = io_inputBit | _GEN_2153; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2155 = i == 10'h272 ? _GEN_2154 : _GEN_2153; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2156 = ~io_inputBit ? 1'h0 : _GEN_2155; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2157 = i == 10'h273 ? _GEN_2156 : _GEN_2155; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2158 = io_inputBit | _GEN_2157; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2159 = i == 10'h273 ? _GEN_2158 : _GEN_2157; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2160 = ~io_inputBit ? 1'h0 : _GEN_2159; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2161 = i == 10'h274 ? _GEN_2160 : _GEN_2159; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2162 = io_inputBit | _GEN_2161; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2163 = i == 10'h274 ? _GEN_2162 : _GEN_2161; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2164 = ~io_inputBit ? 1'h0 : _GEN_2163; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2165 = i == 10'h275 ? _GEN_2164 : _GEN_2163; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2166 = io_inputBit | _GEN_2165; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2167 = i == 10'h275 ? _GEN_2166 : _GEN_2165; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2168 = ~io_inputBit ? 1'h0 : _GEN_2167; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2169 = i == 10'h276 ? _GEN_2168 : _GEN_2167; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2170 = io_inputBit | _GEN_2169; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2171 = i == 10'h276 ? _GEN_2170 : _GEN_2169; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2172 = ~io_inputBit ? 1'h0 : _GEN_2171; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2173 = i == 10'h277 ? _GEN_2172 : _GEN_2171; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2174 = io_inputBit | _GEN_2173; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2175 = i == 10'h277 ? _GEN_2174 : _GEN_2173; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2176 = ~io_inputBit ? 1'h0 : _GEN_2175; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2177 = i == 10'h278 ? _GEN_2176 : _GEN_2175; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2178 = io_inputBit | _GEN_2177; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2179 = i == 10'h278 ? _GEN_2178 : _GEN_2177; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2180 = ~io_inputBit ? 1'h0 : _GEN_2179; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2181 = i == 10'h279 ? _GEN_2180 : _GEN_2179; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2182 = io_inputBit | _GEN_2181; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2183 = i == 10'h279 ? _GEN_2182 : _GEN_2181; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2184 = ~io_inputBit ? 1'h0 : _GEN_2183; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2185 = i == 10'h27a ? _GEN_2184 : _GEN_2183; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2186 = io_inputBit | _GEN_2185; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2187 = i == 10'h27a ? _GEN_2186 : _GEN_2185; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2188 = ~io_inputBit ? 1'h0 : _GEN_2187; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2189 = i == 10'h27b ? _GEN_2188 : _GEN_2187; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2190 = io_inputBit | _GEN_2189; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2191 = i == 10'h27b ? _GEN_2190 : _GEN_2189; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2192 = ~io_inputBit ? 1'h0 : _GEN_2191; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2193 = i == 10'h27c ? _GEN_2192 : _GEN_2191; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2194 = io_inputBit | _GEN_2193; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2195 = i == 10'h27c ? _GEN_2194 : _GEN_2193; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2196 = ~io_inputBit ? 1'h0 : _GEN_2195; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2197 = i == 10'h27d ? _GEN_2196 : _GEN_2195; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2198 = io_inputBit | _GEN_2197; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2199 = i == 10'h27d ? _GEN_2198 : _GEN_2197; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2200 = ~io_inputBit ? 1'h0 : _GEN_2199; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2201 = i == 10'h27e ? _GEN_2200 : _GEN_2199; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2202 = io_inputBit | _GEN_2201; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2203 = i == 10'h27e ? _GEN_2202 : _GEN_2201; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2204 = ~io_inputBit ? 1'h0 : _GEN_2203; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2205 = i == 10'h27f ? _GEN_2204 : _GEN_2203; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2206 = io_inputBit | _GEN_2205; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2207 = i == 10'h27f ? _GEN_2206 : _GEN_2205; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2208 = ~io_inputBit ? 1'h0 : _GEN_2207; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2209 = i == 10'h280 ? _GEN_2208 : _GEN_2207; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2210 = io_inputBit | _GEN_2209; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2211 = i == 10'h280 ? _GEN_2210 : _GEN_2209; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2212 = ~io_inputBit ? 1'h0 : _GEN_2211; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2213 = i == 10'h281 ? _GEN_2212 : _GEN_2211; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2214 = io_inputBit | _GEN_2213; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2215 = i == 10'h281 ? _GEN_2214 : _GEN_2213; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2216 = ~io_inputBit ? 1'h0 : _GEN_2215; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2217 = i == 10'h282 ? _GEN_2216 : _GEN_2215; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2218 = io_inputBit | _GEN_2217; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2219 = i == 10'h282 ? _GEN_2218 : _GEN_2217; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2220 = ~io_inputBit ? 1'h0 : _GEN_2219; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2221 = i == 10'h283 ? _GEN_2220 : _GEN_2219; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2222 = io_inputBit | _GEN_2221; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2223 = i == 10'h283 ? _GEN_2222 : _GEN_2221; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2224 = ~io_inputBit ? 1'h0 : _GEN_2223; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2225 = i == 10'h284 ? _GEN_2224 : _GEN_2223; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2226 = io_inputBit | _GEN_2225; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2227 = i == 10'h284 ? _GEN_2226 : _GEN_2225; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2228 = ~io_inputBit ? 1'h0 : _GEN_2227; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2229 = i == 10'h285 ? _GEN_2228 : _GEN_2227; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2230 = io_inputBit | _GEN_2229; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2231 = i == 10'h285 ? _GEN_2230 : _GEN_2229; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2232 = ~io_inputBit ? 1'h0 : _GEN_2231; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2233 = i == 10'h286 ? _GEN_2232 : _GEN_2231; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2234 = io_inputBit | _GEN_2233; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2235 = i == 10'h286 ? _GEN_2234 : _GEN_2233; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2236 = ~io_inputBit ? 1'h0 : _GEN_2235; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2237 = i == 10'h287 ? _GEN_2236 : _GEN_2235; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2238 = io_inputBit | _GEN_2237; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2239 = i == 10'h287 ? _GEN_2238 : _GEN_2237; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2240 = ~io_inputBit ? 1'h0 : _GEN_2239; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2241 = i == 10'h288 ? _GEN_2240 : _GEN_2239; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2242 = io_inputBit | _GEN_2241; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2243 = i == 10'h288 ? _GEN_2242 : _GEN_2241; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2244 = ~io_inputBit ? 1'h0 : _GEN_2243; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2245 = i == 10'h289 ? _GEN_2244 : _GEN_2243; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2246 = io_inputBit | _GEN_2245; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2247 = i == 10'h289 ? _GEN_2246 : _GEN_2245; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2248 = ~io_inputBit ? 1'h0 : _GEN_2247; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2249 = i == 10'h28a ? _GEN_2248 : _GEN_2247; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2250 = io_inputBit | _GEN_2249; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2251 = i == 10'h28a ? _GEN_2250 : _GEN_2249; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2252 = ~io_inputBit ? 1'h0 : _GEN_2251; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2253 = i == 10'h28b ? _GEN_2252 : _GEN_2251; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2254 = io_inputBit | _GEN_2253; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2255 = i == 10'h28b ? _GEN_2254 : _GEN_2253; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2256 = ~io_inputBit ? 1'h0 : _GEN_2255; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2257 = i == 10'h28c ? _GEN_2256 : _GEN_2255; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2258 = io_inputBit | _GEN_2257; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2259 = i == 10'h28c ? _GEN_2258 : _GEN_2257; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2260 = ~io_inputBit ? 1'h0 : _GEN_2259; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2261 = i == 10'h28d ? _GEN_2260 : _GEN_2259; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2262 = io_inputBit | _GEN_2261; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2263 = i == 10'h28d ? _GEN_2262 : _GEN_2261; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2264 = ~io_inputBit ? 1'h0 : _GEN_2263; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2265 = i == 10'h28e ? _GEN_2264 : _GEN_2263; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2266 = io_inputBit | _GEN_2265; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2267 = i == 10'h28e ? _GEN_2266 : _GEN_2265; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2268 = ~io_inputBit ? 1'h0 : _GEN_2267; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2269 = i == 10'h28f ? _GEN_2268 : _GEN_2267; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2270 = io_inputBit | _GEN_2269; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2271 = i == 10'h28f ? _GEN_2270 : _GEN_2269; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2272 = ~io_inputBit ? 1'h0 : _GEN_2271; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2273 = i == 10'h290 ? _GEN_2272 : _GEN_2271; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2274 = io_inputBit | _GEN_2273; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2275 = i == 10'h290 ? _GEN_2274 : _GEN_2273; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2276 = ~io_inputBit ? 1'h0 : _GEN_2275; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2277 = i == 10'h291 ? _GEN_2276 : _GEN_2275; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2278 = io_inputBit | _GEN_2277; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2279 = i == 10'h291 ? _GEN_2278 : _GEN_2277; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2280 = ~io_inputBit ? 1'h0 : _GEN_2279; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2281 = i == 10'h292 ? _GEN_2280 : _GEN_2279; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2282 = io_inputBit | _GEN_2281; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2283 = i == 10'h292 ? _GEN_2282 : _GEN_2281; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2284 = ~io_inputBit ? 1'h0 : _GEN_2283; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2285 = i == 10'h293 ? _GEN_2284 : _GEN_2283; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2286 = io_inputBit | _GEN_2285; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2287 = i == 10'h293 ? _GEN_2286 : _GEN_2285; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2288 = ~io_inputBit ? 1'h0 : _GEN_2287; // @[lut_mem_online.scala 249:46 251:32]
  wire  _GEN_2289 = i == 10'h294 ? _GEN_2288 : _GEN_2287; // @[lut_mem_online.scala 247:34]
  wire  _GEN_2290 = io_inputBit | _GEN_2289; // @[lut_mem_online.scala 249:46 251:32]
  wire  _T_2295 = counter < 5'h11; // @[lut_mem_online.scala 262:22]
  wire  _T_2297 = counter >= 5'ha; // @[lut_mem_online.scala 270:30]
  wire [4:0] _outResult_T_1 = counter - 5'ha; // @[lut_mem_online.scala 272:41]
  wire  _GEN_2300 = 4'h1 == _outResult_T_1[3:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2301 = 4'h2 == _outResult_T_1[3:0] ? buffer_2 : _GEN_2300; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2302 = 4'h3 == _outResult_T_1[3:0] ? buffer_3 : _GEN_2301; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2303 = 4'h4 == _outResult_T_1[3:0] ? buffer_4 : _GEN_2302; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2304 = 4'h5 == _outResult_T_1[3:0] ? buffer_5 : _GEN_2303; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2305 = 4'h6 == _outResult_T_1[3:0] ? buffer_6 : _GEN_2304; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2306 = 4'h7 == _outResult_T_1[3:0] ? 1'h0 : _GEN_2305; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2307 = 4'h8 == _outResult_T_1[3:0] ? 1'h0 : _GEN_2306; // @[lut_mem_online.scala 272:{23,23}]
  wire  _GEN_2308 = 4'h9 == _outResult_T_1[3:0] ? 1'h0 : _GEN_2307; // @[lut_mem_online.scala 272:{23,23}]
  wire  _T_2301 = ~reset; // @[lut_mem_online.scala 278:21]
  wire  _GEN_2310 = counter >= 5'ha ? _GEN_2308 : outResult; // @[lut_mem_online.scala 270:42 272:23 224:26]
  wire  _GEN_2312 = _T_2 ? 1'h0 : _GEN_2310; // @[lut_mem_online.scala 267:35 269:23]
  wire  _T_2302 = i < 10'h1ff; // @[lut_mem_online.scala 293:18]
  wire [11:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 307:24]
  wire [11:0] _i_T_2 = _i_T + 12'h1; // @[lut_mem_online.scala 307:28]
  wire [11:0] _i_T_5 = _i_T + 12'h2; // @[lut_mem_online.scala 309:28]
  wire [11:0] _GEN_2313 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 308:45 309:17 215:18]
  wire [11:0] _GEN_2314 = _T_10 ? _i_T_2 : _GEN_2313; // @[lut_mem_online.scala 306:39 307:17]
  wire  _T_2307 = i < 10'h3ff; // @[lut_mem_online.scala 316:24]
  wire [9:0] _GEN_2315 = i < 10'h3ff ? 10'h3ff : i; // @[lut_mem_online.scala 316:63 324:15 215:18]
  wire [11:0] _GEN_2316 = i < 10'h1ff ? _GEN_2314 : {{2'd0}, _GEN_2315}; // @[lut_mem_online.scala 293:61]
  wire [4:0] _counter_T_1 = counter + 5'h1; // @[lut_mem_online.scala 327:30]
  wire  _GEN_2318 = counter < 5'h11 & _GEN_2312; // @[lut_mem_online.scala 262:52 335:21]
  wire [11:0] _GEN_2319 = counter < 5'h11 ? _GEN_2316 : {{2'd0}, i}; // @[lut_mem_online.scala 215:18 262:52]
  wire  _GEN_2342 = io_start & _GEN_2318; // @[lut_mem_online.scala 229:29 362:15]
  wire [11:0] _GEN_2343 = io_start ? _GEN_2319 : 12'h0; // @[lut_mem_online.scala 229:29 360:7]
  wire [11:0] _GEN_2346 = reset ? 12'h0 : _GEN_2343; // @[lut_mem_online.scala 215:{18,18}]
  wire  _GEN_2347 = io_start & _T_2295; // @[lut_mem_online.scala 278:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 369:16]
  always @(posedge clock) begin
    i <= _GEN_2346[9:0]; // @[lut_mem_online.scala 215:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h275) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_0 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_0 <= _GEN_883;
          end
        end else begin
          buffer_0 <= _GEN_883;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h285) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_1 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_1 <= _GEN_961;
          end
        end else begin
          buffer_1 <= _GEN_961;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h28d) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_2 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_2 <= _GEN_1081;
          end
        end else begin
          buffer_2 <= _GEN_1081;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h291) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_3 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_3 <= _GEN_1271;
          end
        end else begin
          buffer_3 <= _GEN_1271;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h293) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_4 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_4 <= _GEN_1543;
          end
        end else begin
          buffer_4 <= _GEN_1543;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h294) begin // @[lut_mem_online.scala 247:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 249:46]
            buffer_5 <= 1'h0; // @[lut_mem_online.scala 251:32]
          end else begin
            buffer_5 <= _GEN_1865;
          end
        end else begin
          buffer_5 <= _GEN_1865;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 241:36]
        if (i == 10'h294) begin // @[lut_mem_online.scala 247:34]
          buffer_6 <= _GEN_2290;
        end else if (i == 10'h294) begin // @[lut_mem_online.scala 247:34]
          buffer_6 <= _GEN_2288;
        end else begin
          buffer_6 <= _GEN_2287;
        end
      end
    end
    if (reset) begin // @[lut_mem_online.scala 221:24]
      counter <= 5'h0; // @[lut_mem_online.scala 221:24]
    end else if (io_start) begin // @[lut_mem_online.scala 229:29]
      if (counter < 5'h11) begin // @[lut_mem_online.scala 262:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 327:19]
      end
    end else begin
      counter <= 5'h0; // @[lut_mem_online.scala 361:13]
    end
    if (reset) begin // @[lut_mem_online.scala 224:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 224:26]
    end else begin
      outResult <= _GEN_2342;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_2295 & ~_T_2 & _T_2297 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 278:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2347 & _T_2302 & _T_2301) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 300:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2347 & ~_T_2302 & _T_2307 & _T_2301) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 319:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
