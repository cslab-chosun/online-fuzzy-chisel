module LutMembershipFunctionOnline_4(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [9:0] i; // @[lut_mem_online.scala 206:18]
  reg  buffer_0; // @[lut_mem_online.scala 210:19]
  reg  buffer_1; // @[lut_mem_online.scala 210:19]
  reg  buffer_2; // @[lut_mem_online.scala 210:19]
  reg  buffer_3; // @[lut_mem_online.scala 210:19]
  reg  buffer_4; // @[lut_mem_online.scala 210:19]
  reg  buffer_5; // @[lut_mem_online.scala 210:19]
  reg  buffer_6; // @[lut_mem_online.scala 210:19]
  reg [4:0] counter; // @[lut_mem_online.scala 212:24]
  reg  outResult; // @[lut_mem_online.scala 215:26]
  wire  _T_2 = counter < 5'ha; // @[lut_mem_online.scala 232:22]
  wire  _GEN_0 = i == 10'h0 ? 1'h0 : buffer_0; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_1 = i == 10'h1 ? 1'h0 : _GEN_0; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2 = i == 10'h3 ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_4 = i == 10'h10 ? 1'h0 : i == 10'h7 | _GEN_2; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_6 = i == 10'h44 ? 1'h0 : i == 10'h21 | _GEN_4; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_10 = i == 10'h22a ? 1'h0 : i == 10'h22a | (i == 10'h114 | (i == 10'h89 | _GEN_6)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_11 = i == 10'h0 ? 1'h0 : buffer_1; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_12 = i == 10'h1 ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_13 = i == 10'h3 ? 1'h0 : _GEN_12; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_16 = i == 10'h21 ? 1'h0 : i == 10'h20 | (i == 10'hf | _GEN_13); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_18 = i == 10'h42 ? 1'h0 : i == 10'h22 | _GEN_16; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_20 = i == 10'h46 ? 1'h0 : i == 10'h44 | _GEN_18; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_22 = i == 10'h89 ? 1'h0 : i == 10'h85 | _GEN_20; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_25 = i == 10'h114 ? 1'h0 : i == 10'h10c | (i == 10'h8d | _GEN_22); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_28 = i == 10'h21a ? 1'h0 : i == 10'h21a | (i == 10'h11c | _GEN_25); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_29 = i == 10'h22a ? 1'h0 : _GEN_28; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_32 = i == 10'h23a ? 1'h0 : i == 10'h23a | (i == 10'h22a | _GEN_29); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_33 = i == 10'h0 ? 1'h0 : buffer_2; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_34 = i == 10'h1 ? 1'h0 : _GEN_33; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_35 = i == 10'h8 ? 1'h0 : _GEN_34; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_36 = i == 10'hf ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_37 = i == 10'h11 ? 1'h0 : _GEN_36; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_38 = i == 10'h20 ? 1'h0 : _GEN_37; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_39 = i == 10'h23 ? 1'h0 : _GEN_38; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_41 = i == 10'h43 ? 1'h0 : i == 10'h42 | _GEN_39; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_43 = i == 10'h45 ? 1'h0 : i == 10'h44 | _GEN_41; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_45 = i == 10'h47 ? 1'h0 : i == 10'h46 | _GEN_43; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_46 = i == 10'h85 ? 1'h0 : _GEN_45; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_48 = i == 10'h89 ? 1'h0 : i == 10'h87 | _GEN_46; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_50 = i == 10'h8d ? 1'h0 : i == 10'h8b | _GEN_48; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_52 = i == 10'h10c ? 1'h0 : i == 10'h8f | _GEN_50; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_54 = i == 10'h114 ? 1'h0 : i == 10'h110 | _GEN_52; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_56 = i == 10'h11c ? 1'h0 : i == 10'h118 | _GEN_54; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_58 = i == 10'h21a ? 1'h0 : i == 10'h120 | _GEN_56; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_61 = i == 10'h222 ? 1'h0 : i == 10'h222 | (i == 10'h21a | _GEN_58); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_62 = i == 10'h22a ? 1'h0 : _GEN_61; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_65 = i == 10'h232 ? 1'h0 : i == 10'h232 | (i == 10'h22a | _GEN_62); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_66 = i == 10'h23a ? 1'h0 : _GEN_65; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_69 = i == 10'h242 ? 1'h0 : i == 10'h242 | (i == 10'h23a | _GEN_66); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_70 = i == 10'h0 ? 1'h0 : buffer_3; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_71 = i == 10'h1 ? 1'h0 : _GEN_70; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_72 = i == 10'h8 ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_73 = i == 10'hf ? 1'h0 : _GEN_72; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_74 = i == 10'h11 ? 1'h0 : _GEN_73; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_75 = i == 10'h20 ? 1'h0 : _GEN_74; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_76 = i == 10'h23 ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_77 = i == 10'h85 ? 1'h0 : _GEN_76; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_79 = i == 10'h87 ? 1'h0 : i == 10'h86 | _GEN_77; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_81 = i == 10'h89 ? 1'h0 : i == 10'h88 | _GEN_79; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_83 = i == 10'h8b ? 1'h0 : i == 10'h8a | _GEN_81; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_85 = i == 10'h8d ? 1'h0 : i == 10'h8c | _GEN_83; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_87 = i == 10'h8f ? 1'h0 : i == 10'h8e | _GEN_85; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_89 = i == 10'h10c ? 1'h0 : i == 10'h90 | _GEN_87; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_91 = i == 10'h110 ? 1'h0 : i == 10'h10e | _GEN_89; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_93 = i == 10'h114 ? 1'h0 : i == 10'h112 | _GEN_91; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_95 = i == 10'h118 ? 1'h0 : i == 10'h116 | _GEN_93; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_97 = i == 10'h11c ? 1'h0 : i == 10'h11a | _GEN_95; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_99 = i == 10'h120 ? 1'h0 : i == 10'h11e | _GEN_97; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_101 = i == 10'h21a ? 1'h0 : i == 10'h122 | _GEN_99; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_104 = i == 10'h21e ? 1'h0 : i == 10'h21e | (i == 10'h21a | _GEN_101); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_105 = i == 10'h222 ? 1'h0 : _GEN_104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_108 = i == 10'h226 ? 1'h0 : i == 10'h226 | (i == 10'h222 | _GEN_105); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_109 = i == 10'h22a ? 1'h0 : _GEN_108; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_112 = i == 10'h22e ? 1'h0 : i == 10'h22e | (i == 10'h22a | _GEN_109); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_113 = i == 10'h232 ? 1'h0 : _GEN_112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_116 = i == 10'h236 ? 1'h0 : i == 10'h236 | (i == 10'h232 | _GEN_113); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_117 = i == 10'h23a ? 1'h0 : _GEN_116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_120 = i == 10'h23e ? 1'h0 : i == 10'h23e | (i == 10'h23a | _GEN_117); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_121 = i == 10'h242 ? 1'h0 : _GEN_120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_124 = i == 10'h246 ? 1'h0 : i == 10'h246 | (i == 10'h242 | _GEN_121); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_125 = i == 10'h0 ? 1'h0 : buffer_4; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_126 = i == 10'h1 ? 1'h0 : _GEN_125; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_127 = i == 10'h8 ? 1'h0 : _GEN_126; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_129 = i == 10'h11 ? 1'h0 : i == 10'hf | _GEN_127; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_131 = i == 10'h48 ? 1'h0 : i == 10'h20 | _GEN_129; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_132 = i == 10'h91 ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_134 = i == 10'h10c ? 1'h0 : i == 10'h10b | _GEN_132; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_136 = i == 10'h10e ? 1'h0 : i == 10'h10d | _GEN_134; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_138 = i == 10'h110 ? 1'h0 : i == 10'h10f | _GEN_136; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_140 = i == 10'h112 ? 1'h0 : i == 10'h111 | _GEN_138; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_142 = i == 10'h114 ? 1'h0 : i == 10'h113 | _GEN_140; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_144 = i == 10'h116 ? 1'h0 : i == 10'h115 | _GEN_142; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_146 = i == 10'h118 ? 1'h0 : i == 10'h117 | _GEN_144; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_148 = i == 10'h11a ? 1'h0 : i == 10'h119 | _GEN_146; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_150 = i == 10'h11c ? 1'h0 : i == 10'h11b | _GEN_148; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_152 = i == 10'h11e ? 1'h0 : i == 10'h11d | _GEN_150; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_154 = i == 10'h120 ? 1'h0 : i == 10'h11f | _GEN_152; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_156 = i == 10'h122 ? 1'h0 : i == 10'h121 | _GEN_154; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_159 = i == 10'h218 ? 1'h0 : i == 10'h218 | (i == 10'h123 | _GEN_156); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_160 = i == 10'h21a ? 1'h0 : _GEN_159; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_163 = i == 10'h21c ? 1'h0 : i == 10'h21c | (i == 10'h21a | _GEN_160); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_164 = i == 10'h21e ? 1'h0 : _GEN_163; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_167 = i == 10'h220 ? 1'h0 : i == 10'h220 | (i == 10'h21e | _GEN_164); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_168 = i == 10'h222 ? 1'h0 : _GEN_167; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_171 = i == 10'h224 ? 1'h0 : i == 10'h224 | (i == 10'h222 | _GEN_168); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_172 = i == 10'h226 ? 1'h0 : _GEN_171; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_175 = i == 10'h228 ? 1'h0 : i == 10'h228 | (i == 10'h226 | _GEN_172); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_176 = i == 10'h22a ? 1'h0 : _GEN_175; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_179 = i == 10'h22c ? 1'h0 : i == 10'h22c | (i == 10'h22a | _GEN_176); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_180 = i == 10'h22e ? 1'h0 : _GEN_179; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_183 = i == 10'h230 ? 1'h0 : i == 10'h230 | (i == 10'h22e | _GEN_180); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_184 = i == 10'h232 ? 1'h0 : _GEN_183; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_187 = i == 10'h234 ? 1'h0 : i == 10'h234 | (i == 10'h232 | _GEN_184); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_188 = i == 10'h236 ? 1'h0 : _GEN_187; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_191 = i == 10'h238 ? 1'h0 : i == 10'h238 | (i == 10'h236 | _GEN_188); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_192 = i == 10'h23a ? 1'h0 : _GEN_191; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_195 = i == 10'h23c ? 1'h0 : i == 10'h23c | (i == 10'h23a | _GEN_192); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_196 = i == 10'h23e ? 1'h0 : _GEN_195; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_199 = i == 10'h240 ? 1'h0 : i == 10'h240 | (i == 10'h23e | _GEN_196); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_200 = i == 10'h242 ? 1'h0 : _GEN_199; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_203 = i == 10'h244 ? 1'h0 : i == 10'h244 | (i == 10'h242 | _GEN_200); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_204 = i == 10'h246 ? 1'h0 : _GEN_203; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_207 = i == 10'h248 ? 1'h0 : i == 10'h248 | (i == 10'h246 | _GEN_204); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_208 = i == 10'h0 ? 1'h0 : buffer_5; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_209 = i == 10'h1 ? 1'h0 : _GEN_208; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_210 = i == 10'h8 ? 1'h0 : _GEN_209; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_211 = i == 10'hf ? 1'h0 : _GEN_210; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_212 = i == 10'h11 ? 1'h0 : _GEN_211; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_213 = i == 10'h20 ? 1'h0 : _GEN_212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_214 = i == 10'h48 ? 1'h0 : _GEN_213; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_215 = i == 10'h10b ? 1'h0 : _GEN_214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_216 = i == 10'h124 ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_217 = i == 10'h218 ? 1'h0 : _GEN_216; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_220 = i == 10'h219 ? 1'h0 : i == 10'h219 | (i == 10'h218 | _GEN_217); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_221 = i == 10'h21a ? 1'h0 : _GEN_220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_224 = i == 10'h21b ? 1'h0 : i == 10'h21b | (i == 10'h21a | _GEN_221); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_225 = i == 10'h21c ? 1'h0 : _GEN_224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_228 = i == 10'h21d ? 1'h0 : i == 10'h21d | (i == 10'h21c | _GEN_225); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_229 = i == 10'h21e ? 1'h0 : _GEN_228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_232 = i == 10'h21f ? 1'h0 : i == 10'h21f | (i == 10'h21e | _GEN_229); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_233 = i == 10'h220 ? 1'h0 : _GEN_232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_236 = i == 10'h221 ? 1'h0 : i == 10'h221 | (i == 10'h220 | _GEN_233); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_237 = i == 10'h222 ? 1'h0 : _GEN_236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_240 = i == 10'h223 ? 1'h0 : i == 10'h223 | (i == 10'h222 | _GEN_237); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_241 = i == 10'h224 ? 1'h0 : _GEN_240; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_244 = i == 10'h225 ? 1'h0 : i == 10'h225 | (i == 10'h224 | _GEN_241); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_245 = i == 10'h226 ? 1'h0 : _GEN_244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_248 = i == 10'h227 ? 1'h0 : i == 10'h227 | (i == 10'h226 | _GEN_245); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_249 = i == 10'h228 ? 1'h0 : _GEN_248; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_252 = i == 10'h229 ? 1'h0 : i == 10'h229 | (i == 10'h228 | _GEN_249); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_253 = i == 10'h22a ? 1'h0 : _GEN_252; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_256 = i == 10'h22b ? 1'h0 : i == 10'h22b | (i == 10'h22a | _GEN_253); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_257 = i == 10'h22c ? 1'h0 : _GEN_256; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_260 = i == 10'h22d ? 1'h0 : i == 10'h22d | (i == 10'h22c | _GEN_257); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_261 = i == 10'h22e ? 1'h0 : _GEN_260; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_264 = i == 10'h22f ? 1'h0 : i == 10'h22f | (i == 10'h22e | _GEN_261); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_265 = i == 10'h230 ? 1'h0 : _GEN_264; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_268 = i == 10'h231 ? 1'h0 : i == 10'h231 | (i == 10'h230 | _GEN_265); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_269 = i == 10'h232 ? 1'h0 : _GEN_268; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_272 = i == 10'h233 ? 1'h0 : i == 10'h233 | (i == 10'h232 | _GEN_269); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_273 = i == 10'h234 ? 1'h0 : _GEN_272; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_276 = i == 10'h235 ? 1'h0 : i == 10'h235 | (i == 10'h234 | _GEN_273); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_277 = i == 10'h236 ? 1'h0 : _GEN_276; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_280 = i == 10'h237 ? 1'h0 : i == 10'h237 | (i == 10'h236 | _GEN_277); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_281 = i == 10'h238 ? 1'h0 : _GEN_280; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_284 = i == 10'h239 ? 1'h0 : i == 10'h239 | (i == 10'h238 | _GEN_281); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_285 = i == 10'h23a ? 1'h0 : _GEN_284; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_288 = i == 10'h23b ? 1'h0 : i == 10'h23b | (i == 10'h23a | _GEN_285); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_289 = i == 10'h23c ? 1'h0 : _GEN_288; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_292 = i == 10'h23d ? 1'h0 : i == 10'h23d | (i == 10'h23c | _GEN_289); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_293 = i == 10'h23e ? 1'h0 : _GEN_292; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_296 = i == 10'h23f ? 1'h0 : i == 10'h23f | (i == 10'h23e | _GEN_293); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_297 = i == 10'h240 ? 1'h0 : _GEN_296; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_300 = i == 10'h241 ? 1'h0 : i == 10'h241 | (i == 10'h240 | _GEN_297); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_301 = i == 10'h242 ? 1'h0 : _GEN_300; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_304 = i == 10'h243 ? 1'h0 : i == 10'h243 | (i == 10'h242 | _GEN_301); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_305 = i == 10'h244 ? 1'h0 : _GEN_304; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_308 = i == 10'h245 ? 1'h0 : i == 10'h245 | (i == 10'h244 | _GEN_305); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_309 = i == 10'h246 ? 1'h0 : _GEN_308; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_312 = i == 10'h247 ? 1'h0 : i == 10'h247 | (i == 10'h246 | _GEN_309); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_313 = i == 10'h248 ? 1'h0 : _GEN_312; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_316 = i == 10'h249 ? 1'h0 : i == 10'h249 | (i == 10'h248 | _GEN_313); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_317 = i == 10'h0 ? 1'h0 : buffer_6; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_318 = i == 10'h1 ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_319 = i == 10'h8 ? 1'h0 : _GEN_318; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_320 = i == 10'hf ? 1'h0 : _GEN_319; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_321 = i == 10'h11 ? 1'h0 : _GEN_320; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_322 = i == 10'h20 ? 1'h0 : _GEN_321; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_323 = i == 10'h48 ? 1'h0 : _GEN_322; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_324 = i == 10'h10b ? 1'h0 : _GEN_323; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_325 = i == 10'h124 ? 1'h0 : _GEN_324; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_326 = i == 10'h218 ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_328 = i == 10'h219 ? 1'h0 : i == 10'h218 | _GEN_326; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_330 = i == 10'h21a ? 1'h0 : i == 10'h219 | _GEN_328; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_332 = i == 10'h21b ? 1'h0 : i == 10'h21a | _GEN_330; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_334 = i == 10'h21c ? 1'h0 : i == 10'h21b | _GEN_332; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_336 = i == 10'h21d ? 1'h0 : i == 10'h21c | _GEN_334; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_338 = i == 10'h21e ? 1'h0 : i == 10'h21d | _GEN_336; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_340 = i == 10'h21f ? 1'h0 : i == 10'h21e | _GEN_338; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_342 = i == 10'h220 ? 1'h0 : i == 10'h21f | _GEN_340; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_344 = i == 10'h221 ? 1'h0 : i == 10'h220 | _GEN_342; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_346 = i == 10'h222 ? 1'h0 : i == 10'h221 | _GEN_344; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_348 = i == 10'h223 ? 1'h0 : i == 10'h222 | _GEN_346; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_350 = i == 10'h224 ? 1'h0 : i == 10'h223 | _GEN_348; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_352 = i == 10'h225 ? 1'h0 : i == 10'h224 | _GEN_350; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_354 = i == 10'h226 ? 1'h0 : i == 10'h225 | _GEN_352; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_356 = i == 10'h227 ? 1'h0 : i == 10'h226 | _GEN_354; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_358 = i == 10'h228 ? 1'h0 : i == 10'h227 | _GEN_356; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_360 = i == 10'h229 ? 1'h0 : i == 10'h228 | _GEN_358; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_362 = i == 10'h22a ? 1'h0 : i == 10'h229 | _GEN_360; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_364 = i == 10'h22b ? 1'h0 : i == 10'h22a | _GEN_362; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_366 = i == 10'h22c ? 1'h0 : i == 10'h22b | _GEN_364; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_368 = i == 10'h22d ? 1'h0 : i == 10'h22c | _GEN_366; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_370 = i == 10'h22e ? 1'h0 : i == 10'h22d | _GEN_368; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_372 = i == 10'h22f ? 1'h0 : i == 10'h22e | _GEN_370; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_374 = i == 10'h230 ? 1'h0 : i == 10'h22f | _GEN_372; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_376 = i == 10'h231 ? 1'h0 : i == 10'h230 | _GEN_374; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_378 = i == 10'h232 ? 1'h0 : i == 10'h231 | _GEN_376; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_380 = i == 10'h233 ? 1'h0 : i == 10'h232 | _GEN_378; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_382 = i == 10'h234 ? 1'h0 : i == 10'h233 | _GEN_380; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_384 = i == 10'h235 ? 1'h0 : i == 10'h234 | _GEN_382; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_386 = i == 10'h236 ? 1'h0 : i == 10'h235 | _GEN_384; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_388 = i == 10'h237 ? 1'h0 : i == 10'h236 | _GEN_386; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_390 = i == 10'h238 ? 1'h0 : i == 10'h237 | _GEN_388; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_392 = i == 10'h239 ? 1'h0 : i == 10'h238 | _GEN_390; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_394 = i == 10'h23a ? 1'h0 : i == 10'h239 | _GEN_392; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_396 = i == 10'h23b ? 1'h0 : i == 10'h23a | _GEN_394; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_398 = i == 10'h23c ? 1'h0 : i == 10'h23b | _GEN_396; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_400 = i == 10'h23d ? 1'h0 : i == 10'h23c | _GEN_398; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_402 = i == 10'h23e ? 1'h0 : i == 10'h23d | _GEN_400; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_404 = i == 10'h23f ? 1'h0 : i == 10'h23e | _GEN_402; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_406 = i == 10'h240 ? 1'h0 : i == 10'h23f | _GEN_404; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_408 = i == 10'h241 ? 1'h0 : i == 10'h240 | _GEN_406; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_410 = i == 10'h242 ? 1'h0 : i == 10'h241 | _GEN_408; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_412 = i == 10'h243 ? 1'h0 : i == 10'h242 | _GEN_410; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_414 = i == 10'h244 ? 1'h0 : i == 10'h243 | _GEN_412; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_416 = i == 10'h245 ? 1'h0 : i == 10'h244 | _GEN_414; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_418 = i == 10'h246 ? 1'h0 : i == 10'h245 | _GEN_416; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_420 = i == 10'h247 ? 1'h0 : i == 10'h246 | _GEN_418; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_422 = i == 10'h248 ? 1'h0 : i == 10'h247 | _GEN_420; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_424 = i == 10'h249 ? 1'h0 : i == 10'h248 | _GEN_422; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_426 = i == 10'h0 ? 1'h0 : _GEN_10; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_427 = i == 10'h1 ? 1'h0 : _GEN_426; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_428 = i == 10'h7 ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_430 = i == 10'h10 ? 1'h0 : i == 10'h8 | _GEN_428; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_432 = i == 10'h22 ? 1'h0 : i == 10'h12 | _GEN_430; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_433 = i == 10'h26 ? 1'h0 : _GEN_432; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_438 = i == 10'h11b ? 1'h0 : i == 10'h9c | (i == 10'h8d | (i == 10'h4d | (i == 10'h46 | _GEN_433))); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_440 = i == 10'h13a ? 1'h0 : i == 10'h11b | _GEN_438; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_442 = i == 10'h275 ? 1'h0 : i == 10'h275 | _GEN_440; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_443 = i == 10'h0 ? 1'h0 : _GEN_32; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_444 = i == 10'h4 ? 1'h0 : _GEN_443; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_445 = i == 10'h7 ? 1'h0 : _GEN_444; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_446 = i == 10'h9 ? 1'h0 : _GEN_445; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_448 = i == 10'h13 ? 1'h0 : i == 10'h11 | _GEN_446; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_449 = i == 10'h21 ? 1'h0 : _GEN_448; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_451 = i == 10'h23 ? 1'h0 : i == 10'h22 | _GEN_449; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_452 = i == 10'h25 ? 1'h0 : _GEN_451; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_454 = i == 10'h27 ? 1'h0 : i == 10'h26 | _GEN_452; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_456 = i == 10'h46 ? 1'h0 : i == 10'h44 | _GEN_454; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_459 = i == 10'h4d ? 1'h0 : i == 10'h4b | (i == 10'h48 | _GEN_456); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_462 = i == 10'h8d ? 1'h0 : i == 10'h89 | (i == 10'h4f | _GEN_459); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_465 = i == 10'h9c ? 1'h0 : i == 10'h98 | (i == 10'h91 | _GEN_462); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_467 = i == 10'h113 ? 1'h0 : i == 10'ha0 | _GEN_465; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_470 = i == 10'h11b ? 1'h0 : i == 10'h11b | (i == 10'h113 | _GEN_467); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_471 = i == 10'h123 ? 1'h0 : _GEN_470; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_473 = i == 10'h132 ? 1'h0 : i == 10'h123 | _GEN_471; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_475 = i == 10'h142 ? 1'h0 : i == 10'h13a | _GEN_473; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_477 = i == 10'h265 ? 1'h0 : i == 10'h265 | _GEN_475; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_478 = i == 10'h275 ? 1'h0 : _GEN_477; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_481 = i == 10'h285 ? 1'h0 : i == 10'h285 | (i == 10'h275 | _GEN_478); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_482 = i == 10'h0 ? 1'h0 : _GEN_69; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_483 = i == 10'h4 ? 1'h0 : _GEN_482; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_484 = i == 10'h7 ? 1'h0 : _GEN_483; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_485 = i == 10'h9 ? 1'h0 : _GEN_484; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_486 = i == 10'h11 ? 1'h0 : _GEN_485; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_487 = i == 10'h13 ? 1'h0 : _GEN_486; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_489 = i == 10'h44 ? 1'h0 : i == 10'h43 | _GEN_487; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_491 = i == 10'h46 ? 1'h0 : i == 10'h45 | _GEN_489; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_493 = i == 10'h48 ? 1'h0 : i == 10'h47 | _GEN_491; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_494 = i == 10'h4b ? 1'h0 : _GEN_493; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_496 = i == 10'h4d ? 1'h0 : i == 10'h4c | _GEN_494; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_498 = i == 10'h4f ? 1'h0 : i == 10'h4e | _GEN_496; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_501 = i == 10'h89 ? 1'h0 : i == 10'h87 | (i == 10'h50 | _GEN_498); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_503 = i == 10'h8d ? 1'h0 : i == 10'h8b | _GEN_501; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_505 = i == 10'h91 ? 1'h0 : i == 10'h8f | _GEN_503; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_506 = i == 10'h98 ? 1'h0 : _GEN_505; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_508 = i == 10'h9c ? 1'h0 : i == 10'h9a | _GEN_506; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_510 = i == 10'ha0 ? 1'h0 : i == 10'h9e | _GEN_508; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_512 = i == 10'h10f ? 1'h0 : i == 10'ha2 | _GEN_510; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_515 = i == 10'h113 ? 1'h0 : i == 10'h113 | (i == 10'h10f | _GEN_512); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_516 = i == 10'h117 ? 1'h0 : _GEN_515; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_519 = i == 10'h11b ? 1'h0 : i == 10'h11b | (i == 10'h117 | _GEN_516); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_520 = i == 10'h11f ? 1'h0 : _GEN_519; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_523 = i == 10'h123 ? 1'h0 : i == 10'h123 | (i == 10'h11f | _GEN_520); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_525 = i == 10'h136 ? 1'h0 : i == 10'h132 | _GEN_523; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_527 = i == 10'h13e ? 1'h0 : i == 10'h13a | _GEN_525; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_529 = i == 10'h146 ? 1'h0 : i == 10'h142 | _GEN_527; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_530 = i == 10'h265 ? 1'h0 : _GEN_529; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_533 = i == 10'h26d ? 1'h0 : i == 10'h26d | (i == 10'h265 | _GEN_530); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_534 = i == 10'h275 ? 1'h0 : _GEN_533; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_537 = i == 10'h27d ? 1'h0 : i == 10'h27d | (i == 10'h275 | _GEN_534); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_538 = i == 10'h285 ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_541 = i == 10'h28d ? 1'h0 : i == 10'h28d | (i == 10'h285 | _GEN_538); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_542 = i == 10'h0 ? 1'h0 : _GEN_124; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_543 = i == 10'h4 ? 1'h0 : _GEN_542; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_544 = i == 10'h9 ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_545 = i == 10'hf ? 1'h0 : _GEN_544; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_546 = i == 10'h11 ? 1'h0 : _GEN_545; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_547 = i == 10'h20 ? 1'h0 : _GEN_546; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_548 = i == 10'h28 ? 1'h0 : _GEN_547; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_549 = i == 10'h42 ? 1'h0 : _GEN_548; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_550 = i == 10'h48 ? 1'h0 : _GEN_549; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_551 = i == 10'h4b ? 1'h0 : _GEN_550; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_552 = i == 10'h51 ? 1'h0 : _GEN_551; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_554 = i == 10'h87 ? 1'h0 : i == 10'h86 | _GEN_552; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_556 = i == 10'h89 ? 1'h0 : i == 10'h88 | _GEN_554; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_558 = i == 10'h8b ? 1'h0 : i == 10'h8a | _GEN_556; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_560 = i == 10'h8d ? 1'h0 : i == 10'h8c | _GEN_558; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_562 = i == 10'h8f ? 1'h0 : i == 10'h8e | _GEN_560; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_564 = i == 10'h91 ? 1'h0 : i == 10'h90 | _GEN_562; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_565 = i == 10'h98 ? 1'h0 : _GEN_564; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_567 = i == 10'h9a ? 1'h0 : i == 10'h99 | _GEN_565; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_569 = i == 10'h9c ? 1'h0 : i == 10'h9b | _GEN_567; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_571 = i == 10'h9e ? 1'h0 : i == 10'h9d | _GEN_569; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_573 = i == 10'ha0 ? 1'h0 : i == 10'h9f | _GEN_571; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_575 = i == 10'ha2 ? 1'h0 : i == 10'ha1 | _GEN_573; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_577 = i == 10'h10d ? 1'h0 : i == 10'ha3 | _GEN_575; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_580 = i == 10'h10f ? 1'h0 : i == 10'h10f | (i == 10'h10d | _GEN_577); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_581 = i == 10'h111 ? 1'h0 : _GEN_580; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_584 = i == 10'h113 ? 1'h0 : i == 10'h113 | (i == 10'h111 | _GEN_581); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_585 = i == 10'h115 ? 1'h0 : _GEN_584; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_588 = i == 10'h117 ? 1'h0 : i == 10'h117 | (i == 10'h115 | _GEN_585); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_589 = i == 10'h119 ? 1'h0 : _GEN_588; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_592 = i == 10'h11b ? 1'h0 : i == 10'h11b | (i == 10'h119 | _GEN_589); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_593 = i == 10'h11d ? 1'h0 : _GEN_592; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_596 = i == 10'h11f ? 1'h0 : i == 10'h11f | (i == 10'h11d | _GEN_593); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_597 = i == 10'h121 ? 1'h0 : _GEN_596; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_600 = i == 10'h123 ? 1'h0 : i == 10'h123 | (i == 10'h121 | _GEN_597); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_602 = i == 10'h134 ? 1'h0 : i == 10'h132 | _GEN_600; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_604 = i == 10'h138 ? 1'h0 : i == 10'h136 | _GEN_602; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_606 = i == 10'h13c ? 1'h0 : i == 10'h13a | _GEN_604; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_608 = i == 10'h140 ? 1'h0 : i == 10'h13e | _GEN_606; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_610 = i == 10'h144 ? 1'h0 : i == 10'h142 | _GEN_608; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_612 = i == 10'h148 ? 1'h0 : i == 10'h146 | _GEN_610; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_613 = i == 10'h265 ? 1'h0 : _GEN_612; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_616 = i == 10'h269 ? 1'h0 : i == 10'h269 | (i == 10'h265 | _GEN_613); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_617 = i == 10'h26d ? 1'h0 : _GEN_616; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_620 = i == 10'h271 ? 1'h0 : i == 10'h271 | (i == 10'h26d | _GEN_617); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_621 = i == 10'h275 ? 1'h0 : _GEN_620; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_624 = i == 10'h279 ? 1'h0 : i == 10'h279 | (i == 10'h275 | _GEN_621); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_625 = i == 10'h27d ? 1'h0 : _GEN_624; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_628 = i == 10'h281 ? 1'h0 : i == 10'h281 | (i == 10'h27d | _GEN_625); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_629 = i == 10'h285 ? 1'h0 : _GEN_628; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_632 = i == 10'h289 ? 1'h0 : i == 10'h289 | (i == 10'h285 | _GEN_629); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_633 = i == 10'h28d ? 1'h0 : _GEN_632; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_636 = i == 10'h291 ? 1'h0 : i == 10'h291 | (i == 10'h28d | _GEN_633); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_637 = i == 10'h0 ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_638 = i == 10'h4 ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_639 = i == 10'h9 ? 1'h0 : _GEN_638; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_640 = i == 10'hf ? 1'h0 : _GEN_639; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_642 = i == 10'h20 ? 1'h0 : i == 10'h11 | _GEN_640; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_643 = i == 10'h28 ? 1'h0 : _GEN_642; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_646 = i == 10'h85 ? 1'h0 : i == 10'h4b | (i == 10'h48 | _GEN_643); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_647 = i == 10'ha4 ? 1'h0 : _GEN_646; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_648 = i == 10'h10c ? 1'h0 : _GEN_647; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_651 = i == 10'h10d ? 1'h0 : i == 10'h10d | (i == 10'h10c | _GEN_648); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_652 = i == 10'h10e ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_655 = i == 10'h10f ? 1'h0 : i == 10'h10f | (i == 10'h10e | _GEN_652); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_656 = i == 10'h110 ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_659 = i == 10'h111 ? 1'h0 : i == 10'h111 | (i == 10'h110 | _GEN_656); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_660 = i == 10'h112 ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_663 = i == 10'h113 ? 1'h0 : i == 10'h113 | (i == 10'h112 | _GEN_660); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_664 = i == 10'h114 ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_667 = i == 10'h115 ? 1'h0 : i == 10'h115 | (i == 10'h114 | _GEN_664); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_668 = i == 10'h116 ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_671 = i == 10'h117 ? 1'h0 : i == 10'h117 | (i == 10'h116 | _GEN_668); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_672 = i == 10'h118 ? 1'h0 : _GEN_671; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_675 = i == 10'h119 ? 1'h0 : i == 10'h119 | (i == 10'h118 | _GEN_672); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_676 = i == 10'h11a ? 1'h0 : _GEN_675; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_679 = i == 10'h11b ? 1'h0 : i == 10'h11b | (i == 10'h11a | _GEN_676); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_680 = i == 10'h11c ? 1'h0 : _GEN_679; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_683 = i == 10'h11d ? 1'h0 : i == 10'h11d | (i == 10'h11c | _GEN_680); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_684 = i == 10'h11e ? 1'h0 : _GEN_683; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_687 = i == 10'h11f ? 1'h0 : i == 10'h11f | (i == 10'h11e | _GEN_684); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_688 = i == 10'h120 ? 1'h0 : _GEN_687; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_691 = i == 10'h121 ? 1'h0 : i == 10'h121 | (i == 10'h120 | _GEN_688); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_692 = i == 10'h122 ? 1'h0 : _GEN_691; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_695 = i == 10'h123 ? 1'h0 : i == 10'h123 | (i == 10'h122 | _GEN_692); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_696 = i == 10'h124 ? 1'h0 : _GEN_695; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_698 = i == 10'h131 ? 1'h0 : i == 10'h124 | _GEN_696; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_700 = i == 10'h133 ? 1'h0 : i == 10'h132 | _GEN_698; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_702 = i == 10'h135 ? 1'h0 : i == 10'h134 | _GEN_700; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_704 = i == 10'h137 ? 1'h0 : i == 10'h136 | _GEN_702; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_706 = i == 10'h139 ? 1'h0 : i == 10'h138 | _GEN_704; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_708 = i == 10'h13b ? 1'h0 : i == 10'h13a | _GEN_706; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_710 = i == 10'h13d ? 1'h0 : i == 10'h13c | _GEN_708; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_712 = i == 10'h13f ? 1'h0 : i == 10'h13e | _GEN_710; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_714 = i == 10'h141 ? 1'h0 : i == 10'h140 | _GEN_712; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_716 = i == 10'h143 ? 1'h0 : i == 10'h142 | _GEN_714; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_718 = i == 10'h145 ? 1'h0 : i == 10'h144 | _GEN_716; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_720 = i == 10'h147 ? 1'h0 : i == 10'h146 | _GEN_718; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_722 = i == 10'h149 ? 1'h0 : i == 10'h148 | _GEN_720; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_724 = i == 10'h263 ? 1'h0 : i == 10'h263 | _GEN_722; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_725 = i == 10'h265 ? 1'h0 : _GEN_724; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_728 = i == 10'h267 ? 1'h0 : i == 10'h267 | (i == 10'h265 | _GEN_725); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_729 = i == 10'h269 ? 1'h0 : _GEN_728; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_732 = i == 10'h26b ? 1'h0 : i == 10'h26b | (i == 10'h269 | _GEN_729); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_733 = i == 10'h26d ? 1'h0 : _GEN_732; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_736 = i == 10'h26f ? 1'h0 : i == 10'h26f | (i == 10'h26d | _GEN_733); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_737 = i == 10'h271 ? 1'h0 : _GEN_736; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_740 = i == 10'h273 ? 1'h0 : i == 10'h273 | (i == 10'h271 | _GEN_737); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_741 = i == 10'h275 ? 1'h0 : _GEN_740; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_744 = i == 10'h277 ? 1'h0 : i == 10'h277 | (i == 10'h275 | _GEN_741); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_745 = i == 10'h279 ? 1'h0 : _GEN_744; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_748 = i == 10'h27b ? 1'h0 : i == 10'h27b | (i == 10'h279 | _GEN_745); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_749 = i == 10'h27d ? 1'h0 : _GEN_748; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_752 = i == 10'h27f ? 1'h0 : i == 10'h27f | (i == 10'h27d | _GEN_749); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_753 = i == 10'h281 ? 1'h0 : _GEN_752; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_756 = i == 10'h283 ? 1'h0 : i == 10'h283 | (i == 10'h281 | _GEN_753); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_757 = i == 10'h285 ? 1'h0 : _GEN_756; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_760 = i == 10'h287 ? 1'h0 : i == 10'h287 | (i == 10'h285 | _GEN_757); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_761 = i == 10'h289 ? 1'h0 : _GEN_760; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_764 = i == 10'h28b ? 1'h0 : i == 10'h28b | (i == 10'h289 | _GEN_761); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_765 = i == 10'h28d ? 1'h0 : _GEN_764; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_768 = i == 10'h28f ? 1'h0 : i == 10'h28f | (i == 10'h28d | _GEN_765); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_769 = i == 10'h291 ? 1'h0 : _GEN_768; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_772 = i == 10'h293 ? 1'h0 : i == 10'h293 | (i == 10'h291 | _GEN_769); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_773 = i == 10'h0 ? 1'h0 : _GEN_316; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_774 = i == 10'h4 ? 1'h0 : _GEN_773; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_775 = i == 10'h9 ? 1'h0 : _GEN_774; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_776 = i == 10'hf ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_777 = i == 10'h11 ? 1'h0 : _GEN_776; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_778 = i == 10'h20 ? 1'h0 : _GEN_777; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_779 = i == 10'h28 ? 1'h0 : _GEN_778; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_780 = i == 10'h48 ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_781 = i == 10'h4b ? 1'h0 : _GEN_780; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_782 = i == 10'h85 ? 1'h0 : _GEN_781; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_783 = i == 10'ha4 ? 1'h0 : _GEN_782; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_785 = i == 10'h10c ? 1'h0 : i == 10'h10c | _GEN_783; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_787 = i == 10'h10d ? 1'h0 : i == 10'h10d | _GEN_785; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_789 = i == 10'h10e ? 1'h0 : i == 10'h10e | _GEN_787; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_791 = i == 10'h10f ? 1'h0 : i == 10'h10f | _GEN_789; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_793 = i == 10'h110 ? 1'h0 : i == 10'h110 | _GEN_791; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_795 = i == 10'h111 ? 1'h0 : i == 10'h111 | _GEN_793; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_797 = i == 10'h112 ? 1'h0 : i == 10'h112 | _GEN_795; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_799 = i == 10'h113 ? 1'h0 : i == 10'h113 | _GEN_797; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_801 = i == 10'h114 ? 1'h0 : i == 10'h114 | _GEN_799; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_803 = i == 10'h115 ? 1'h0 : i == 10'h115 | _GEN_801; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_805 = i == 10'h116 ? 1'h0 : i == 10'h116 | _GEN_803; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_807 = i == 10'h117 ? 1'h0 : i == 10'h117 | _GEN_805; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_809 = i == 10'h118 ? 1'h0 : i == 10'h118 | _GEN_807; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_811 = i == 10'h119 ? 1'h0 : i == 10'h119 | _GEN_809; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_813 = i == 10'h11a ? 1'h0 : i == 10'h11a | _GEN_811; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_815 = i == 10'h11b ? 1'h0 : i == 10'h11b | _GEN_813; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_817 = i == 10'h11c ? 1'h0 : i == 10'h11c | _GEN_815; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_819 = i == 10'h11d ? 1'h0 : i == 10'h11d | _GEN_817; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_821 = i == 10'h11e ? 1'h0 : i == 10'h11e | _GEN_819; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_823 = i == 10'h11f ? 1'h0 : i == 10'h11f | _GEN_821; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_825 = i == 10'h120 ? 1'h0 : i == 10'h120 | _GEN_823; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_827 = i == 10'h121 ? 1'h0 : i == 10'h121 | _GEN_825; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_829 = i == 10'h122 ? 1'h0 : i == 10'h122 | _GEN_827; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_831 = i == 10'h123 ? 1'h0 : i == 10'h123 | _GEN_829; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_833 = i == 10'h124 ? 1'h0 : i == 10'h124 | _GEN_831; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_834 = i == 10'h263 ? 1'h0 : _GEN_833; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_837 = i == 10'h264 ? 1'h0 : i == 10'h264 | (i == 10'h263 | _GEN_834); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_838 = i == 10'h265 ? 1'h0 : _GEN_837; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_841 = i == 10'h266 ? 1'h0 : i == 10'h266 | (i == 10'h265 | _GEN_838); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_842 = i == 10'h267 ? 1'h0 : _GEN_841; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_845 = i == 10'h268 ? 1'h0 : i == 10'h268 | (i == 10'h267 | _GEN_842); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_846 = i == 10'h269 ? 1'h0 : _GEN_845; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_849 = i == 10'h26a ? 1'h0 : i == 10'h26a | (i == 10'h269 | _GEN_846); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_850 = i == 10'h26b ? 1'h0 : _GEN_849; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_853 = i == 10'h26c ? 1'h0 : i == 10'h26c | (i == 10'h26b | _GEN_850); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_854 = i == 10'h26d ? 1'h0 : _GEN_853; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_857 = i == 10'h26e ? 1'h0 : i == 10'h26e | (i == 10'h26d | _GEN_854); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_858 = i == 10'h26f ? 1'h0 : _GEN_857; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_861 = i == 10'h270 ? 1'h0 : i == 10'h270 | (i == 10'h26f | _GEN_858); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_862 = i == 10'h271 ? 1'h0 : _GEN_861; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_865 = i == 10'h272 ? 1'h0 : i == 10'h272 | (i == 10'h271 | _GEN_862); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_866 = i == 10'h273 ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_869 = i == 10'h274 ? 1'h0 : i == 10'h274 | (i == 10'h273 | _GEN_866); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_870 = i == 10'h275 ? 1'h0 : _GEN_869; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_873 = i == 10'h276 ? 1'h0 : i == 10'h276 | (i == 10'h275 | _GEN_870); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_874 = i == 10'h277 ? 1'h0 : _GEN_873; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_877 = i == 10'h278 ? 1'h0 : i == 10'h278 | (i == 10'h277 | _GEN_874); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_878 = i == 10'h279 ? 1'h0 : _GEN_877; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_881 = i == 10'h27a ? 1'h0 : i == 10'h27a | (i == 10'h279 | _GEN_878); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_882 = i == 10'h27b ? 1'h0 : _GEN_881; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_885 = i == 10'h27c ? 1'h0 : i == 10'h27c | (i == 10'h27b | _GEN_882); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_886 = i == 10'h27d ? 1'h0 : _GEN_885; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_889 = i == 10'h27e ? 1'h0 : i == 10'h27e | (i == 10'h27d | _GEN_886); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_890 = i == 10'h27f ? 1'h0 : _GEN_889; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_893 = i == 10'h280 ? 1'h0 : i == 10'h280 | (i == 10'h27f | _GEN_890); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_894 = i == 10'h281 ? 1'h0 : _GEN_893; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_897 = i == 10'h282 ? 1'h0 : i == 10'h282 | (i == 10'h281 | _GEN_894); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_898 = i == 10'h283 ? 1'h0 : _GEN_897; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_901 = i == 10'h284 ? 1'h0 : i == 10'h284 | (i == 10'h283 | _GEN_898); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_902 = i == 10'h285 ? 1'h0 : _GEN_901; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_905 = i == 10'h286 ? 1'h0 : i == 10'h286 | (i == 10'h285 | _GEN_902); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_906 = i == 10'h287 ? 1'h0 : _GEN_905; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_909 = i == 10'h288 ? 1'h0 : i == 10'h288 | (i == 10'h287 | _GEN_906); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_910 = i == 10'h289 ? 1'h0 : _GEN_909; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_913 = i == 10'h28a ? 1'h0 : i == 10'h28a | (i == 10'h289 | _GEN_910); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_914 = i == 10'h28b ? 1'h0 : _GEN_913; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_917 = i == 10'h28c ? 1'h0 : i == 10'h28c | (i == 10'h28b | _GEN_914); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_918 = i == 10'h28d ? 1'h0 : _GEN_917; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_921 = i == 10'h28e ? 1'h0 : i == 10'h28e | (i == 10'h28d | _GEN_918); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_922 = i == 10'h28f ? 1'h0 : _GEN_921; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_925 = i == 10'h290 ? 1'h0 : i == 10'h290 | (i == 10'h28f | _GEN_922); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_926 = i == 10'h291 ? 1'h0 : _GEN_925; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_929 = i == 10'h292 ? 1'h0 : i == 10'h292 | (i == 10'h291 | _GEN_926); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_930 = i == 10'h293 ? 1'h0 : _GEN_929; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_933 = i == 10'h294 ? 1'h0 : i == 10'h294 | (i == 10'h293 | _GEN_930); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_934 = i == 10'h0 ? 1'h0 : i == 10'h249 | _GEN_424; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_935 = i == 10'h4 ? 1'h0 : _GEN_934; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_936 = i == 10'h9 ? 1'h0 : _GEN_935; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_937 = i == 10'hf ? 1'h0 : _GEN_936; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_938 = i == 10'h11 ? 1'h0 : _GEN_937; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_939 = i == 10'h20 ? 1'h0 : _GEN_938; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_940 = i == 10'h28 ? 1'h0 : _GEN_939; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_941 = i == 10'h48 ? 1'h0 : _GEN_940; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_942 = i == 10'h4b ? 1'h0 : _GEN_941; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_943 = i == 10'ha4 ? 1'h0 : _GEN_942; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_944 = i == 10'h10b ? 1'h0 : _GEN_943; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_945 = i == 10'h124 ? 1'h0 : _GEN_944; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_946 = i == 10'h218 ? 1'h0 : _GEN_945; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_948 = i == 10'h219 ? 1'h0 : i == 10'h218 | _GEN_946; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_950 = i == 10'h21a ? 1'h0 : i == 10'h219 | _GEN_948; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_952 = i == 10'h21b ? 1'h0 : i == 10'h21a | _GEN_950; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_954 = i == 10'h21c ? 1'h0 : i == 10'h21b | _GEN_952; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_956 = i == 10'h21d ? 1'h0 : i == 10'h21c | _GEN_954; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_958 = i == 10'h21e ? 1'h0 : i == 10'h21d | _GEN_956; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_960 = i == 10'h21f ? 1'h0 : i == 10'h21e | _GEN_958; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_962 = i == 10'h220 ? 1'h0 : i == 10'h21f | _GEN_960; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_964 = i == 10'h221 ? 1'h0 : i == 10'h220 | _GEN_962; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_966 = i == 10'h222 ? 1'h0 : i == 10'h221 | _GEN_964; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_968 = i == 10'h223 ? 1'h0 : i == 10'h222 | _GEN_966; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_970 = i == 10'h224 ? 1'h0 : i == 10'h223 | _GEN_968; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_972 = i == 10'h225 ? 1'h0 : i == 10'h224 | _GEN_970; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_974 = i == 10'h226 ? 1'h0 : i == 10'h225 | _GEN_972; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_976 = i == 10'h227 ? 1'h0 : i == 10'h226 | _GEN_974; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_978 = i == 10'h228 ? 1'h0 : i == 10'h227 | _GEN_976; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_980 = i == 10'h229 ? 1'h0 : i == 10'h228 | _GEN_978; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_982 = i == 10'h22a ? 1'h0 : i == 10'h229 | _GEN_980; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_984 = i == 10'h22b ? 1'h0 : i == 10'h22a | _GEN_982; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_986 = i == 10'h22c ? 1'h0 : i == 10'h22b | _GEN_984; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_988 = i == 10'h22d ? 1'h0 : i == 10'h22c | _GEN_986; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_990 = i == 10'h22e ? 1'h0 : i == 10'h22d | _GEN_988; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_992 = i == 10'h22f ? 1'h0 : i == 10'h22e | _GEN_990; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_994 = i == 10'h230 ? 1'h0 : i == 10'h22f | _GEN_992; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_996 = i == 10'h231 ? 1'h0 : i == 10'h230 | _GEN_994; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_998 = i == 10'h232 ? 1'h0 : i == 10'h231 | _GEN_996; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1000 = i == 10'h233 ? 1'h0 : i == 10'h232 | _GEN_998; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1002 = i == 10'h234 ? 1'h0 : i == 10'h233 | _GEN_1000; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1004 = i == 10'h235 ? 1'h0 : i == 10'h234 | _GEN_1002; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1006 = i == 10'h236 ? 1'h0 : i == 10'h235 | _GEN_1004; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1008 = i == 10'h237 ? 1'h0 : i == 10'h236 | _GEN_1006; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1010 = i == 10'h238 ? 1'h0 : i == 10'h237 | _GEN_1008; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1012 = i == 10'h239 ? 1'h0 : i == 10'h238 | _GEN_1010; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1014 = i == 10'h23a ? 1'h0 : i == 10'h239 | _GEN_1012; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1016 = i == 10'h23b ? 1'h0 : i == 10'h23a | _GEN_1014; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1018 = i == 10'h23c ? 1'h0 : i == 10'h23b | _GEN_1016; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1020 = i == 10'h23d ? 1'h0 : i == 10'h23c | _GEN_1018; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1022 = i == 10'h23e ? 1'h0 : i == 10'h23d | _GEN_1020; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1024 = i == 10'h23f ? 1'h0 : i == 10'h23e | _GEN_1022; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1026 = i == 10'h240 ? 1'h0 : i == 10'h23f | _GEN_1024; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1028 = i == 10'h241 ? 1'h0 : i == 10'h240 | _GEN_1026; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1030 = i == 10'h242 ? 1'h0 : i == 10'h241 | _GEN_1028; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1032 = i == 10'h243 ? 1'h0 : i == 10'h242 | _GEN_1030; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1034 = i == 10'h244 ? 1'h0 : i == 10'h243 | _GEN_1032; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1036 = i == 10'h245 ? 1'h0 : i == 10'h244 | _GEN_1034; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1038 = i == 10'h246 ? 1'h0 : i == 10'h245 | _GEN_1036; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1040 = i == 10'h247 ? 1'h0 : i == 10'h246 | _GEN_1038; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1042 = i == 10'h248 ? 1'h0 : i == 10'h247 | _GEN_1040; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1044 = i == 10'h249 ? 1'h0 : i == 10'h248 | _GEN_1042; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1046 = i == 10'h263 ? 1'h0 : i == 10'h249 | _GEN_1044; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1048 = i == 10'h264 ? 1'h0 : i == 10'h263 | _GEN_1046; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1050 = i == 10'h265 ? 1'h0 : i == 10'h264 | _GEN_1048; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1052 = i == 10'h266 ? 1'h0 : i == 10'h265 | _GEN_1050; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1054 = i == 10'h267 ? 1'h0 : i == 10'h266 | _GEN_1052; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1056 = i == 10'h268 ? 1'h0 : i == 10'h267 | _GEN_1054; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1058 = i == 10'h269 ? 1'h0 : i == 10'h268 | _GEN_1056; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1060 = i == 10'h26a ? 1'h0 : i == 10'h269 | _GEN_1058; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1062 = i == 10'h26b ? 1'h0 : i == 10'h26a | _GEN_1060; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1064 = i == 10'h26c ? 1'h0 : i == 10'h26b | _GEN_1062; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1066 = i == 10'h26d ? 1'h0 : i == 10'h26c | _GEN_1064; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1068 = i == 10'h26e ? 1'h0 : i == 10'h26d | _GEN_1066; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1070 = i == 10'h26f ? 1'h0 : i == 10'h26e | _GEN_1068; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1072 = i == 10'h270 ? 1'h0 : i == 10'h26f | _GEN_1070; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1074 = i == 10'h271 ? 1'h0 : i == 10'h270 | _GEN_1072; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1076 = i == 10'h272 ? 1'h0 : i == 10'h271 | _GEN_1074; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1078 = i == 10'h273 ? 1'h0 : i == 10'h272 | _GEN_1076; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1080 = i == 10'h274 ? 1'h0 : i == 10'h273 | _GEN_1078; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1082 = i == 10'h275 ? 1'h0 : i == 10'h274 | _GEN_1080; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1084 = i == 10'h276 ? 1'h0 : i == 10'h275 | _GEN_1082; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1086 = i == 10'h277 ? 1'h0 : i == 10'h276 | _GEN_1084; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1088 = i == 10'h278 ? 1'h0 : i == 10'h277 | _GEN_1086; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1090 = i == 10'h279 ? 1'h0 : i == 10'h278 | _GEN_1088; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1092 = i == 10'h27a ? 1'h0 : i == 10'h279 | _GEN_1090; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1094 = i == 10'h27b ? 1'h0 : i == 10'h27a | _GEN_1092; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1096 = i == 10'h27c ? 1'h0 : i == 10'h27b | _GEN_1094; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1098 = i == 10'h27d ? 1'h0 : i == 10'h27c | _GEN_1096; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1100 = i == 10'h27e ? 1'h0 : i == 10'h27d | _GEN_1098; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1102 = i == 10'h27f ? 1'h0 : i == 10'h27e | _GEN_1100; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1104 = i == 10'h280 ? 1'h0 : i == 10'h27f | _GEN_1102; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1106 = i == 10'h281 ? 1'h0 : i == 10'h280 | _GEN_1104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1108 = i == 10'h282 ? 1'h0 : i == 10'h281 | _GEN_1106; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1110 = i == 10'h283 ? 1'h0 : i == 10'h282 | _GEN_1108; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1112 = i == 10'h284 ? 1'h0 : i == 10'h283 | _GEN_1110; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1114 = i == 10'h285 ? 1'h0 : i == 10'h284 | _GEN_1112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1116 = i == 10'h286 ? 1'h0 : i == 10'h285 | _GEN_1114; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1118 = i == 10'h287 ? 1'h0 : i == 10'h286 | _GEN_1116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1120 = i == 10'h288 ? 1'h0 : i == 10'h287 | _GEN_1118; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1122 = i == 10'h289 ? 1'h0 : i == 10'h288 | _GEN_1120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1124 = i == 10'h28a ? 1'h0 : i == 10'h289 | _GEN_1122; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1126 = i == 10'h28b ? 1'h0 : i == 10'h28a | _GEN_1124; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1128 = i == 10'h28c ? 1'h0 : i == 10'h28b | _GEN_1126; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1130 = i == 10'h28d ? 1'h0 : i == 10'h28c | _GEN_1128; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1132 = i == 10'h28e ? 1'h0 : i == 10'h28d | _GEN_1130; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1134 = i == 10'h28f ? 1'h0 : i == 10'h28e | _GEN_1132; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1136 = i == 10'h290 ? 1'h0 : i == 10'h28f | _GEN_1134; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1138 = i == 10'h291 ? 1'h0 : i == 10'h290 | _GEN_1136; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1140 = i == 10'h292 ? 1'h0 : i == 10'h291 | _GEN_1138; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1142 = i == 10'h293 ? 1'h0 : i == 10'h292 | _GEN_1140; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1144 = i == 10'h294 ? 1'h0 : i == 10'h293 | _GEN_1142; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1146 = i == 10'h0 ? 1'h0 : _GEN_442; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1147 = i == 10'h1 ? 1'h0 : _GEN_1146; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1148 = i == 10'h4 ? 1'h0 : _GEN_1147; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1149 = i == 10'h9 ? 1'h0 : _GEN_1148; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1151 = i == 10'h28 ? 1'h0 : i == 10'h27 | _GEN_1149; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1152 = i == 10'h4f ? 1'h0 : _GEN_1151; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1156 = i == 10'h14a ? 1'h0 : i == 10'ha4 | (i == 10'h51 | (i == 10'h4f | _GEN_1152)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1158 = i == 10'h295 ? 1'h0 : i == 10'h295 | _GEN_1156; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1159 = i == 10'h0 ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1160 = i == 10'h3 ? 1'h0 : _GEN_1159; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1161 = i == 10'h4 ? 1'h0 : _GEN_1160; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1162 = i == 10'h8 ? 1'h0 : _GEN_1161; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1163 = i == 10'h9 ? 1'h0 : _GEN_1162; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1164 = i == 10'h12 ? 1'h0 : _GEN_1163; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1166 = i == 10'h27 ? 1'h0 : i == 10'h26 | _GEN_1164; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1167 = i == 10'h28 ? 1'h0 : _GEN_1166; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1168 = i == 10'h4d ? 1'h0 : _GEN_1167; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1171 = i == 10'h4f ? 1'h0 : i == 10'h4f | (i == 10'h4d | _GEN_1168); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1172 = i == 10'h51 ? 1'h0 : _GEN_1171; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1174 = i == 10'h14a ? 1'h0 : i == 10'ha4 | _GEN_1172; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1176 = i == 10'h295 ? 1'h0 : i == 10'h295 | _GEN_1174; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1177 = i == 10'h0 ? 1'h0 : _GEN_541; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1178 = i == 10'h3 ? 1'h0 : _GEN_1177; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1179 = i == 10'h4 ? 1'h0 : _GEN_1178; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1180 = i == 10'h8 ? 1'h0 : _GEN_1179; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1181 = i == 10'h9 ? 1'h0 : _GEN_1180; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1182 = i == 10'h25 ? 1'h0 : _GEN_1181; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1183 = i == 10'h28 ? 1'h0 : _GEN_1182; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1184 = i == 10'h4c ? 1'h0 : _GEN_1183; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1187 = i == 10'h4d ? 1'h0 : i == 10'h4d | (i == 10'h4c | _GEN_1184); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1188 = i == 10'h4e ? 1'h0 : _GEN_1187; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1191 = i == 10'h4f ? 1'h0 : i == 10'h4f | (i == 10'h4e | _GEN_1188); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1192 = i == 10'h50 ? 1'h0 : _GEN_1191; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1195 = i == 10'h51 ? 1'h0 : i == 10'h51 | (i == 10'h50 | _GEN_1192); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1196 = i == 10'h0 ? 1'h0 : _GEN_636; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1197 = i == 10'h3 ? 1'h0 : _GEN_1196; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1198 = i == 10'h4 ? 1'h0 : _GEN_1197; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1199 = i == 10'h8 ? 1'h0 : _GEN_1198; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1200 = i == 10'h9 ? 1'h0 : _GEN_1199; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1201 = i == 10'h25 ? 1'h0 : _GEN_1200; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1202 = i == 10'h28 ? 1'h0 : _GEN_1201; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1204 = i == 10'h4c ? 1'h0 : i == 10'h4c | _GEN_1202; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1206 = i == 10'h4d ? 1'h0 : i == 10'h4d | _GEN_1204; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1208 = i == 10'h4e ? 1'h0 : i == 10'h4e | _GEN_1206; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1210 = i == 10'h4f ? 1'h0 : i == 10'h4f | _GEN_1208; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1212 = i == 10'h50 ? 1'h0 : i == 10'h50 | _GEN_1210; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1214 = i == 10'h51 ? 1'h0 : i == 10'h51 | _GEN_1212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1215 = i == 10'h0 ? 1'h0 : _GEN_772; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1216 = i == 10'h3 ? 1'h0 : _GEN_1215; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1217 = i == 10'h4 ? 1'h0 : _GEN_1216; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1218 = i == 10'h8 ? 1'h0 : _GEN_1217; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1219 = i == 10'h9 ? 1'h0 : _GEN_1218; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1220 = i == 10'h28 ? 1'h0 : _GEN_1219; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1221 = i == 10'h4b ? 1'h0 : _GEN_1220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1222 = i == 10'h98 ? 1'h0 : _GEN_1221; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1224 = i == 10'h99 ? 1'h0 : i == 10'h98 | _GEN_1222; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1226 = i == 10'h9a ? 1'h0 : i == 10'h99 | _GEN_1224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1228 = i == 10'h9b ? 1'h0 : i == 10'h9a | _GEN_1226; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1230 = i == 10'h9c ? 1'h0 : i == 10'h9b | _GEN_1228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1232 = i == 10'h9d ? 1'h0 : i == 10'h9c | _GEN_1230; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1234 = i == 10'h9e ? 1'h0 : i == 10'h9d | _GEN_1232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1236 = i == 10'h9f ? 1'h0 : i == 10'h9e | _GEN_1234; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1238 = i == 10'ha0 ? 1'h0 : i == 10'h9f | _GEN_1236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1240 = i == 10'ha1 ? 1'h0 : i == 10'ha0 | _GEN_1238; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1242 = i == 10'ha2 ? 1'h0 : i == 10'ha1 | _GEN_1240; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1244 = i == 10'ha3 ? 1'h0 : i == 10'ha2 | _GEN_1242; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1246 = i == 10'ha4 ? 1'h0 : i == 10'ha3 | _GEN_1244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1247 = i == 10'h14a ? 1'h0 : _GEN_1246; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1249 = i == 10'h295 ? 1'h0 : i == 10'h295 | _GEN_1247; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1250 = i == 10'h0 ? 1'h0 : _GEN_933; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1251 = i == 10'h3 ? 1'h0 : _GEN_1250; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1252 = i == 10'h4 ? 1'h0 : _GEN_1251; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1253 = i == 10'h8 ? 1'h0 : _GEN_1252; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1254 = i == 10'h9 ? 1'h0 : _GEN_1253; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1255 = i == 10'h28 ? 1'h0 : _GEN_1254; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1256 = i == 10'h4b ? 1'h0 : _GEN_1255; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1257 = i == 10'ha4 ? 1'h0 : _GEN_1256; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1258 = i == 10'h131 ? 1'h0 : _GEN_1257; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1260 = i == 10'h132 ? 1'h0 : i == 10'h131 | _GEN_1258; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1262 = i == 10'h133 ? 1'h0 : i == 10'h132 | _GEN_1260; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1264 = i == 10'h134 ? 1'h0 : i == 10'h133 | _GEN_1262; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1266 = i == 10'h135 ? 1'h0 : i == 10'h134 | _GEN_1264; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1268 = i == 10'h136 ? 1'h0 : i == 10'h135 | _GEN_1266; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1270 = i == 10'h137 ? 1'h0 : i == 10'h136 | _GEN_1268; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1272 = i == 10'h138 ? 1'h0 : i == 10'h137 | _GEN_1270; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1274 = i == 10'h139 ? 1'h0 : i == 10'h138 | _GEN_1272; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1276 = i == 10'h13a ? 1'h0 : i == 10'h139 | _GEN_1274; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1278 = i == 10'h13b ? 1'h0 : i == 10'h13a | _GEN_1276; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1280 = i == 10'h13c ? 1'h0 : i == 10'h13b | _GEN_1278; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1282 = i == 10'h13d ? 1'h0 : i == 10'h13c | _GEN_1280; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1284 = i == 10'h13e ? 1'h0 : i == 10'h13d | _GEN_1282; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1286 = i == 10'h13f ? 1'h0 : i == 10'h13e | _GEN_1284; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1288 = i == 10'h140 ? 1'h0 : i == 10'h13f | _GEN_1286; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1290 = i == 10'h141 ? 1'h0 : i == 10'h140 | _GEN_1288; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1292 = i == 10'h142 ? 1'h0 : i == 10'h141 | _GEN_1290; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1294 = i == 10'h143 ? 1'h0 : i == 10'h142 | _GEN_1292; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1296 = i == 10'h144 ? 1'h0 : i == 10'h143 | _GEN_1294; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1298 = i == 10'h145 ? 1'h0 : i == 10'h144 | _GEN_1296; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1300 = i == 10'h146 ? 1'h0 : i == 10'h145 | _GEN_1298; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1302 = i == 10'h147 ? 1'h0 : i == 10'h146 | _GEN_1300; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1304 = i == 10'h148 ? 1'h0 : i == 10'h147 | _GEN_1302; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1306 = i == 10'h149 ? 1'h0 : i == 10'h148 | _GEN_1304; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1308 = i == 10'h0 ? 1'h0 : i == 10'h294 | _GEN_1144; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1309 = i == 10'h3 ? 1'h0 : _GEN_1308; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1310 = i == 10'h4 ? 1'h0 : _GEN_1309; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1311 = i == 10'h8 ? 1'h0 : _GEN_1310; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1312 = i == 10'h9 ? 1'h0 : _GEN_1311; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1313 = i == 10'h28 ? 1'h0 : _GEN_1312; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1314 = i == 10'h4b ? 1'h0 : _GEN_1313; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1315 = i == 10'ha4 ? 1'h0 : _GEN_1314; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1316 = i == 10'h263 ? 1'h0 : _GEN_1315; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1318 = i == 10'h264 ? 1'h0 : i == 10'h263 | _GEN_1316; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1320 = i == 10'h265 ? 1'h0 : i == 10'h264 | _GEN_1318; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1322 = i == 10'h266 ? 1'h0 : i == 10'h265 | _GEN_1320; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1324 = i == 10'h267 ? 1'h0 : i == 10'h266 | _GEN_1322; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1326 = i == 10'h268 ? 1'h0 : i == 10'h267 | _GEN_1324; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1328 = i == 10'h269 ? 1'h0 : i == 10'h268 | _GEN_1326; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1330 = i == 10'h26a ? 1'h0 : i == 10'h269 | _GEN_1328; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1332 = i == 10'h26b ? 1'h0 : i == 10'h26a | _GEN_1330; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1334 = i == 10'h26c ? 1'h0 : i == 10'h26b | _GEN_1332; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1336 = i == 10'h26d ? 1'h0 : i == 10'h26c | _GEN_1334; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1338 = i == 10'h26e ? 1'h0 : i == 10'h26d | _GEN_1336; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1340 = i == 10'h26f ? 1'h0 : i == 10'h26e | _GEN_1338; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1342 = i == 10'h270 ? 1'h0 : i == 10'h26f | _GEN_1340; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1344 = i == 10'h271 ? 1'h0 : i == 10'h270 | _GEN_1342; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1346 = i == 10'h272 ? 1'h0 : i == 10'h271 | _GEN_1344; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1348 = i == 10'h273 ? 1'h0 : i == 10'h272 | _GEN_1346; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1350 = i == 10'h274 ? 1'h0 : i == 10'h273 | _GEN_1348; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1352 = i == 10'h275 ? 1'h0 : i == 10'h274 | _GEN_1350; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1354 = i == 10'h276 ? 1'h0 : i == 10'h275 | _GEN_1352; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1356 = i == 10'h277 ? 1'h0 : i == 10'h276 | _GEN_1354; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1358 = i == 10'h278 ? 1'h0 : i == 10'h277 | _GEN_1356; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1360 = i == 10'h279 ? 1'h0 : i == 10'h278 | _GEN_1358; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1362 = i == 10'h27a ? 1'h0 : i == 10'h279 | _GEN_1360; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1364 = i == 10'h27b ? 1'h0 : i == 10'h27a | _GEN_1362; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1366 = i == 10'h27c ? 1'h0 : i == 10'h27b | _GEN_1364; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1368 = i == 10'h27d ? 1'h0 : i == 10'h27c | _GEN_1366; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1370 = i == 10'h27e ? 1'h0 : i == 10'h27d | _GEN_1368; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1372 = i == 10'h27f ? 1'h0 : i == 10'h27e | _GEN_1370; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1374 = i == 10'h280 ? 1'h0 : i == 10'h27f | _GEN_1372; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1376 = i == 10'h281 ? 1'h0 : i == 10'h280 | _GEN_1374; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1378 = i == 10'h282 ? 1'h0 : i == 10'h281 | _GEN_1376; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1380 = i == 10'h283 ? 1'h0 : i == 10'h282 | _GEN_1378; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1382 = i == 10'h284 ? 1'h0 : i == 10'h283 | _GEN_1380; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1384 = i == 10'h285 ? 1'h0 : i == 10'h284 | _GEN_1382; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1386 = i == 10'h286 ? 1'h0 : i == 10'h285 | _GEN_1384; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1388 = i == 10'h287 ? 1'h0 : i == 10'h286 | _GEN_1386; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1390 = i == 10'h288 ? 1'h0 : i == 10'h287 | _GEN_1388; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1392 = i == 10'h289 ? 1'h0 : i == 10'h288 | _GEN_1390; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1394 = i == 10'h28a ? 1'h0 : i == 10'h289 | _GEN_1392; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1396 = i == 10'h28b ? 1'h0 : i == 10'h28a | _GEN_1394; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1398 = i == 10'h28c ? 1'h0 : i == 10'h28b | _GEN_1396; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1400 = i == 10'h28d ? 1'h0 : i == 10'h28c | _GEN_1398; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1402 = i == 10'h28e ? 1'h0 : i == 10'h28d | _GEN_1400; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1404 = i == 10'h28f ? 1'h0 : i == 10'h28e | _GEN_1402; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1406 = i == 10'h290 ? 1'h0 : i == 10'h28f | _GEN_1404; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1408 = i == 10'h291 ? 1'h0 : i == 10'h290 | _GEN_1406; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1410 = i == 10'h292 ? 1'h0 : i == 10'h291 | _GEN_1408; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1412 = i == 10'h293 ? 1'h0 : i == 10'h292 | _GEN_1410; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1414 = i == 10'h294 ? 1'h0 : i == 10'h293 | _GEN_1412; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1416 = i == 10'h0 ? 1'h0 : _GEN_1158; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1417 = i == 10'h1 ? 1'h0 : _GEN_1416; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1418 = i == 10'h4 ? 1'h0 : _GEN_1417; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1421 = i == 10'h2b ? 1'h0 : i == 10'h16 | (i == 10'h15 | _GEN_1418); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1422 = i == 10'h2e ? 1'h0 : _GEN_1421; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1423 = i == 10'h58 ? 1'h0 : _GEN_1422; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1424 = i == 10'h5d ? 1'h0 : _GEN_1423; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1425 = i == 10'hb2 ? 1'h0 : _GEN_1424; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1427 = i == 10'h166 ? 1'h0 : i == 10'hbb | _GEN_1425; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1431 = i == 10'h2f2 ? 1'h0 : i == 10'h2f2 | (i == 10'h178 | (i == 10'h166 | _GEN_1427)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1432 = i == 10'h1 ? 1'h0 : _GEN_1176; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1433 = i == 10'h2 ? 1'h0 : _GEN_1432; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1434 = i == 10'h5 ? 1'h0 : _GEN_1433; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1435 = i == 10'h9 ? 1'h0 : _GEN_1434; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1436 = i == 10'hb ? 1'h0 : _GEN_1435; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1437 = i == 10'h14 ? 1'h0 : _GEN_1436; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1438 = i == 10'h17 ? 1'h0 : _GEN_1437; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1439 = i == 10'h2a ? 1'h0 : _GEN_1438; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1441 = i == 10'h2c ? 1'h0 : i == 10'h2b | _GEN_1439; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1442 = i == 10'h2d ? 1'h0 : _GEN_1441; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1444 = i == 10'h2f ? 1'h0 : i == 10'h2e | _GEN_1442; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1445 = i == 10'h56 ? 1'h0 : _GEN_1444; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1447 = i == 10'h5a ? 1'h0 : i == 10'h58 | _GEN_1445; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1448 = i == 10'h5b ? 1'h0 : _GEN_1447; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1450 = i == 10'h5f ? 1'h0 : i == 10'h5d | _GEN_1448; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1451 = i == 10'hae ? 1'h0 : _GEN_1450; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1453 = i == 10'hb6 ? 1'h0 : i == 10'hb2 | _GEN_1451; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1455 = i == 10'hbb ? 1'h0 : i == 10'hb7 | _GEN_1453; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1457 = i == 10'h15e ? 1'h0 : i == 10'hbf | _GEN_1455; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1460 = i == 10'h166 ? 1'h0 : i == 10'h166 | (i == 10'h15e | _GEN_1457); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1461 = i == 10'h16e ? 1'h0 : _GEN_1460; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1464 = i == 10'h178 ? 1'h0 : i == 10'h170 | (i == 10'h16e | _GEN_1461); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1467 = i == 10'h2e2 ? 1'h0 : i == 10'h2e2 | (i == 10'h180 | _GEN_1464); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1468 = i == 10'h2f2 ? 1'h0 : _GEN_1467; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1471 = i == 10'h302 ? 1'h0 : i == 10'h302 | (i == 10'h2f2 | _GEN_1468); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1472 = i == 10'h1 ? 1'h0 : _GEN_1195; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1473 = i == 10'h2 ? 1'h0 : _GEN_1472; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1474 = i == 10'h5 ? 1'h0 : _GEN_1473; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1475 = i == 10'h9 ? 1'h0 : _GEN_1474; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1476 = i == 10'hb ? 1'h0 : _GEN_1475; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1477 = i == 10'h14 ? 1'h0 : _GEN_1476; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1478 = i == 10'h17 ? 1'h0 : _GEN_1477; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1479 = i == 10'h55 ? 1'h0 : _GEN_1478; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1481 = i == 10'h57 ? 1'h0 : i == 10'h56 | _GEN_1479; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1483 = i == 10'h59 ? 1'h0 : i == 10'h58 | _GEN_1481; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1486 = i == 10'h5c ? 1'h0 : i == 10'h5b | (i == 10'h5a | _GEN_1483); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1488 = i == 10'h5e ? 1'h0 : i == 10'h5d | _GEN_1486; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1490 = i == 10'h60 ? 1'h0 : i == 10'h5f | _GEN_1488; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1491 = i == 10'hac ? 1'h0 : _GEN_1490; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1493 = i == 10'hb0 ? 1'h0 : i == 10'hae | _GEN_1491; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1495 = i == 10'hb4 ? 1'h0 : i == 10'hb2 | _GEN_1493; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1497 = i == 10'hb7 ? 1'h0 : i == 10'hb6 | _GEN_1495; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1499 = i == 10'hbb ? 1'h0 : i == 10'hb9 | _GEN_1497; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1501 = i == 10'hbf ? 1'h0 : i == 10'hbd | _GEN_1499; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1503 = i == 10'h15a ? 1'h0 : i == 10'hc1 | _GEN_1501; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1506 = i == 10'h15e ? 1'h0 : i == 10'h15e | (i == 10'h15a | _GEN_1503); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1507 = i == 10'h162 ? 1'h0 : _GEN_1506; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1510 = i == 10'h166 ? 1'h0 : i == 10'h166 | (i == 10'h162 | _GEN_1507); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1511 = i == 10'h16a ? 1'h0 : _GEN_1510; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1514 = i == 10'h16e ? 1'h0 : i == 10'h16e | (i == 10'h16a | _GEN_1511); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1515 = i == 10'h170 ? 1'h0 : _GEN_1514; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1517 = i == 10'h178 ? 1'h0 : i == 10'h174 | _GEN_1515; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1519 = i == 10'h180 ? 1'h0 : i == 10'h17c | _GEN_1517; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1521 = i == 10'h2e2 ? 1'h0 : i == 10'h184 | _GEN_1519; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1524 = i == 10'h2ea ? 1'h0 : i == 10'h2ea | (i == 10'h2e2 | _GEN_1521); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1525 = i == 10'h2f2 ? 1'h0 : _GEN_1524; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1528 = i == 10'h2fa ? 1'h0 : i == 10'h2fa | (i == 10'h2f2 | _GEN_1525); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1529 = i == 10'h302 ? 1'h0 : _GEN_1528; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1532 = i == 10'h30a ? 1'h0 : i == 10'h30a | (i == 10'h302 | _GEN_1529); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1533 = i == 10'h1 ? 1'h0 : _GEN_1214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1534 = i == 10'h2 ? 1'h0 : _GEN_1533; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1535 = i == 10'h5 ? 1'h0 : _GEN_1534; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1536 = i == 10'h9 ? 1'h0 : _GEN_1535; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1537 = i == 10'hb ? 1'h0 : _GEN_1536; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1538 = i == 10'h14 ? 1'h0 : _GEN_1537; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1539 = i == 10'h17 ? 1'h0 : _GEN_1538; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1540 = i == 10'hab ? 1'h0 : _GEN_1539; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1542 = i == 10'had ? 1'h0 : i == 10'hac | _GEN_1540; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1544 = i == 10'haf ? 1'h0 : i == 10'hae | _GEN_1542; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1546 = i == 10'hb1 ? 1'h0 : i == 10'hb0 | _GEN_1544; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1548 = i == 10'hb3 ? 1'h0 : i == 10'hb2 | _GEN_1546; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1550 = i == 10'hb5 ? 1'h0 : i == 10'hb4 | _GEN_1548; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1552 = i == 10'hb7 ? 1'h0 : i == 10'hb6 | _GEN_1550; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1554 = i == 10'hb9 ? 1'h0 : i == 10'hb8 | _GEN_1552; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1556 = i == 10'hbb ? 1'h0 : i == 10'hba | _GEN_1554; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1558 = i == 10'hbd ? 1'h0 : i == 10'hbc | _GEN_1556; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1560 = i == 10'hbf ? 1'h0 : i == 10'hbe | _GEN_1558; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1562 = i == 10'hc1 ? 1'h0 : i == 10'hc0 | _GEN_1560; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1564 = i == 10'h158 ? 1'h0 : i == 10'hc2 | _GEN_1562; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1567 = i == 10'h15a ? 1'h0 : i == 10'h15a | (i == 10'h158 | _GEN_1564); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1568 = i == 10'h15c ? 1'h0 : _GEN_1567; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1571 = i == 10'h15e ? 1'h0 : i == 10'h15e | (i == 10'h15c | _GEN_1568); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1572 = i == 10'h160 ? 1'h0 : _GEN_1571; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1575 = i == 10'h162 ? 1'h0 : i == 10'h162 | (i == 10'h160 | _GEN_1572); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1576 = i == 10'h164 ? 1'h0 : _GEN_1575; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1579 = i == 10'h166 ? 1'h0 : i == 10'h166 | (i == 10'h164 | _GEN_1576); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1580 = i == 10'h168 ? 1'h0 : _GEN_1579; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1583 = i == 10'h16a ? 1'h0 : i == 10'h16a | (i == 10'h168 | _GEN_1580); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1584 = i == 10'h16c ? 1'h0 : _GEN_1583; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1587 = i == 10'h16e ? 1'h0 : i == 10'h16e | (i == 10'h16c | _GEN_1584); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1588 = i == 10'h170 ? 1'h0 : _GEN_1587; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1590 = i == 10'h174 ? 1'h0 : i == 10'h172 | _GEN_1588; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1592 = i == 10'h178 ? 1'h0 : i == 10'h176 | _GEN_1590; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1594 = i == 10'h17c ? 1'h0 : i == 10'h17a | _GEN_1592; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1596 = i == 10'h180 ? 1'h0 : i == 10'h17e | _GEN_1594; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1598 = i == 10'h184 ? 1'h0 : i == 10'h182 | _GEN_1596; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1600 = i == 10'h2e2 ? 1'h0 : i == 10'h186 | _GEN_1598; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1603 = i == 10'h2e6 ? 1'h0 : i == 10'h2e6 | (i == 10'h2e2 | _GEN_1600); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1604 = i == 10'h2ea ? 1'h0 : _GEN_1603; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1607 = i == 10'h2ee ? 1'h0 : i == 10'h2ee | (i == 10'h2ea | _GEN_1604); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1608 = i == 10'h2f2 ? 1'h0 : _GEN_1607; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1611 = i == 10'h2f6 ? 1'h0 : i == 10'h2f6 | (i == 10'h2f2 | _GEN_1608); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1612 = i == 10'h2fa ? 1'h0 : _GEN_1611; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1615 = i == 10'h2fe ? 1'h0 : i == 10'h2fe | (i == 10'h2fa | _GEN_1612); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1616 = i == 10'h302 ? 1'h0 : _GEN_1615; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1619 = i == 10'h306 ? 1'h0 : i == 10'h306 | (i == 10'h302 | _GEN_1616); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1620 = i == 10'h30a ? 1'h0 : _GEN_1619; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1623 = i == 10'h30e ? 1'h0 : i == 10'h30e | (i == 10'h30a | _GEN_1620); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1624 = i == 10'h1 ? 1'h0 : _GEN_1249; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1625 = i == 10'h2 ? 1'h0 : _GEN_1624; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1626 = i == 10'h5 ? 1'h0 : _GEN_1625; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1627 = i == 10'h9 ? 1'h0 : _GEN_1626; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1628 = i == 10'hb ? 1'h0 : _GEN_1627; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1629 = i == 10'h14 ? 1'h0 : _GEN_1628; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1630 = i == 10'h30 ? 1'h0 : _GEN_1629; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1631 = i == 10'h61 ? 1'h0 : _GEN_1630; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1632 = i == 10'hc3 ? 1'h0 : _GEN_1631; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1633 = i == 10'h157 ? 1'h0 : _GEN_1632; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1636 = i == 10'h158 ? 1'h0 : i == 10'h158 | (i == 10'h157 | _GEN_1633); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1637 = i == 10'h159 ? 1'h0 : _GEN_1636; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1640 = i == 10'h15a ? 1'h0 : i == 10'h15a | (i == 10'h159 | _GEN_1637); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1641 = i == 10'h15b ? 1'h0 : _GEN_1640; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1644 = i == 10'h15c ? 1'h0 : i == 10'h15c | (i == 10'h15b | _GEN_1641); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1645 = i == 10'h15d ? 1'h0 : _GEN_1644; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1648 = i == 10'h15e ? 1'h0 : i == 10'h15e | (i == 10'h15d | _GEN_1645); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1649 = i == 10'h15f ? 1'h0 : _GEN_1648; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1652 = i == 10'h160 ? 1'h0 : i == 10'h160 | (i == 10'h15f | _GEN_1649); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1653 = i == 10'h161 ? 1'h0 : _GEN_1652; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1656 = i == 10'h162 ? 1'h0 : i == 10'h162 | (i == 10'h161 | _GEN_1653); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1657 = i == 10'h163 ? 1'h0 : _GEN_1656; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1660 = i == 10'h164 ? 1'h0 : i == 10'h164 | (i == 10'h163 | _GEN_1657); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1661 = i == 10'h165 ? 1'h0 : _GEN_1660; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1664 = i == 10'h166 ? 1'h0 : i == 10'h166 | (i == 10'h165 | _GEN_1661); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1665 = i == 10'h167 ? 1'h0 : _GEN_1664; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1668 = i == 10'h168 ? 1'h0 : i == 10'h168 | (i == 10'h167 | _GEN_1665); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1669 = i == 10'h169 ? 1'h0 : _GEN_1668; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1672 = i == 10'h16a ? 1'h0 : i == 10'h16a | (i == 10'h169 | _GEN_1669); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1673 = i == 10'h16b ? 1'h0 : _GEN_1672; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1676 = i == 10'h16c ? 1'h0 : i == 10'h16c | (i == 10'h16b | _GEN_1673); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1677 = i == 10'h16d ? 1'h0 : _GEN_1676; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1680 = i == 10'h16e ? 1'h0 : i == 10'h16e | (i == 10'h16d | _GEN_1677); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1681 = i == 10'h16f ? 1'h0 : _GEN_1680; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1682 = i == 10'h170 ? 1'h0 : _GEN_1681; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1684 = i == 10'h172 ? 1'h0 : i == 10'h171 | _GEN_1682; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1686 = i == 10'h174 ? 1'h0 : i == 10'h173 | _GEN_1684; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1688 = i == 10'h176 ? 1'h0 : i == 10'h175 | _GEN_1686; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1690 = i == 10'h178 ? 1'h0 : i == 10'h177 | _GEN_1688; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1692 = i == 10'h17a ? 1'h0 : i == 10'h179 | _GEN_1690; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1694 = i == 10'h17c ? 1'h0 : i == 10'h17b | _GEN_1692; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1696 = i == 10'h17e ? 1'h0 : i == 10'h17d | _GEN_1694; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1698 = i == 10'h180 ? 1'h0 : i == 10'h17f | _GEN_1696; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1700 = i == 10'h182 ? 1'h0 : i == 10'h181 | _GEN_1698; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1702 = i == 10'h184 ? 1'h0 : i == 10'h183 | _GEN_1700; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1704 = i == 10'h186 ? 1'h0 : i == 10'h185 | _GEN_1702; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1707 = i == 10'h2e0 ? 1'h0 : i == 10'h2e0 | (i == 10'h187 | _GEN_1704); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1708 = i == 10'h2e2 ? 1'h0 : _GEN_1707; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1711 = i == 10'h2e4 ? 1'h0 : i == 10'h2e4 | (i == 10'h2e2 | _GEN_1708); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1712 = i == 10'h2e6 ? 1'h0 : _GEN_1711; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1715 = i == 10'h2e8 ? 1'h0 : i == 10'h2e8 | (i == 10'h2e6 | _GEN_1712); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1716 = i == 10'h2ea ? 1'h0 : _GEN_1715; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1719 = i == 10'h2ec ? 1'h0 : i == 10'h2ec | (i == 10'h2ea | _GEN_1716); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1720 = i == 10'h2ee ? 1'h0 : _GEN_1719; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1723 = i == 10'h2f0 ? 1'h0 : i == 10'h2f0 | (i == 10'h2ee | _GEN_1720); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1724 = i == 10'h2f2 ? 1'h0 : _GEN_1723; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1727 = i == 10'h2f4 ? 1'h0 : i == 10'h2f4 | (i == 10'h2f2 | _GEN_1724); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1728 = i == 10'h2f6 ? 1'h0 : _GEN_1727; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1731 = i == 10'h2f8 ? 1'h0 : i == 10'h2f8 | (i == 10'h2f6 | _GEN_1728); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1732 = i == 10'h2fa ? 1'h0 : _GEN_1731; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1735 = i == 10'h2fc ? 1'h0 : i == 10'h2fc | (i == 10'h2fa | _GEN_1732); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1736 = i == 10'h2fe ? 1'h0 : _GEN_1735; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1739 = i == 10'h300 ? 1'h0 : i == 10'h300 | (i == 10'h2fe | _GEN_1736); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1740 = i == 10'h302 ? 1'h0 : _GEN_1739; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1743 = i == 10'h304 ? 1'h0 : i == 10'h304 | (i == 10'h302 | _GEN_1740); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1744 = i == 10'h306 ? 1'h0 : _GEN_1743; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1747 = i == 10'h308 ? 1'h0 : i == 10'h308 | (i == 10'h306 | _GEN_1744); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1748 = i == 10'h30a ? 1'h0 : _GEN_1747; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1751 = i == 10'h30c ? 1'h0 : i == 10'h30c | (i == 10'h30a | _GEN_1748); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1752 = i == 10'h30e ? 1'h0 : _GEN_1751; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1755 = i == 10'h310 ? 1'h0 : i == 10'h310 | (i == 10'h30e | _GEN_1752); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1756 = i == 10'h1 ? 1'h0 : i == 10'h149 | _GEN_1306; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1757 = i == 10'h2 ? 1'h0 : _GEN_1756; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1758 = i == 10'h5 ? 1'h0 : _GEN_1757; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1759 = i == 10'h9 ? 1'h0 : _GEN_1758; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1760 = i == 10'hb ? 1'h0 : _GEN_1759; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1761 = i == 10'h14 ? 1'h0 : _GEN_1760; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1762 = i == 10'h30 ? 1'h0 : _GEN_1761; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1763 = i == 10'h61 ? 1'h0 : _GEN_1762; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1765 = i == 10'h157 ? 1'h0 : i == 10'h157 | _GEN_1763; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1767 = i == 10'h158 ? 1'h0 : i == 10'h158 | _GEN_1765; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1769 = i == 10'h159 ? 1'h0 : i == 10'h159 | _GEN_1767; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1771 = i == 10'h15a ? 1'h0 : i == 10'h15a | _GEN_1769; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1773 = i == 10'h15b ? 1'h0 : i == 10'h15b | _GEN_1771; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1775 = i == 10'h15c ? 1'h0 : i == 10'h15c | _GEN_1773; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1777 = i == 10'h15d ? 1'h0 : i == 10'h15d | _GEN_1775; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1779 = i == 10'h15e ? 1'h0 : i == 10'h15e | _GEN_1777; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1781 = i == 10'h15f ? 1'h0 : i == 10'h15f | _GEN_1779; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1783 = i == 10'h160 ? 1'h0 : i == 10'h160 | _GEN_1781; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1785 = i == 10'h161 ? 1'h0 : i == 10'h161 | _GEN_1783; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1787 = i == 10'h162 ? 1'h0 : i == 10'h162 | _GEN_1785; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1789 = i == 10'h163 ? 1'h0 : i == 10'h163 | _GEN_1787; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1791 = i == 10'h164 ? 1'h0 : i == 10'h164 | _GEN_1789; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1793 = i == 10'h165 ? 1'h0 : i == 10'h165 | _GEN_1791; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1795 = i == 10'h166 ? 1'h0 : i == 10'h166 | _GEN_1793; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1797 = i == 10'h167 ? 1'h0 : i == 10'h167 | _GEN_1795; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1799 = i == 10'h168 ? 1'h0 : i == 10'h168 | _GEN_1797; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1801 = i == 10'h169 ? 1'h0 : i == 10'h169 | _GEN_1799; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1803 = i == 10'h16a ? 1'h0 : i == 10'h16a | _GEN_1801; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1805 = i == 10'h16b ? 1'h0 : i == 10'h16b | _GEN_1803; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1807 = i == 10'h16c ? 1'h0 : i == 10'h16c | _GEN_1805; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1809 = i == 10'h16d ? 1'h0 : i == 10'h16d | _GEN_1807; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1811 = i == 10'h16e ? 1'h0 : i == 10'h16e | _GEN_1809; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1813 = i == 10'h188 ? 1'h0 : i == 10'h16f | _GEN_1811; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1814 = i == 10'h2e0 ? 1'h0 : _GEN_1813; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1817 = i == 10'h2e1 ? 1'h0 : i == 10'h2e1 | (i == 10'h2e0 | _GEN_1814); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1818 = i == 10'h2e2 ? 1'h0 : _GEN_1817; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1821 = i == 10'h2e3 ? 1'h0 : i == 10'h2e3 | (i == 10'h2e2 | _GEN_1818); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1822 = i == 10'h2e4 ? 1'h0 : _GEN_1821; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1825 = i == 10'h2e5 ? 1'h0 : i == 10'h2e5 | (i == 10'h2e4 | _GEN_1822); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1826 = i == 10'h2e6 ? 1'h0 : _GEN_1825; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1829 = i == 10'h2e7 ? 1'h0 : i == 10'h2e7 | (i == 10'h2e6 | _GEN_1826); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1830 = i == 10'h2e8 ? 1'h0 : _GEN_1829; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1833 = i == 10'h2e9 ? 1'h0 : i == 10'h2e9 | (i == 10'h2e8 | _GEN_1830); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1834 = i == 10'h2ea ? 1'h0 : _GEN_1833; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1837 = i == 10'h2eb ? 1'h0 : i == 10'h2eb | (i == 10'h2ea | _GEN_1834); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1838 = i == 10'h2ec ? 1'h0 : _GEN_1837; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1841 = i == 10'h2ed ? 1'h0 : i == 10'h2ed | (i == 10'h2ec | _GEN_1838); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1842 = i == 10'h2ee ? 1'h0 : _GEN_1841; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1845 = i == 10'h2ef ? 1'h0 : i == 10'h2ef | (i == 10'h2ee | _GEN_1842); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1846 = i == 10'h2f0 ? 1'h0 : _GEN_1845; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1849 = i == 10'h2f1 ? 1'h0 : i == 10'h2f1 | (i == 10'h2f0 | _GEN_1846); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1850 = i == 10'h2f2 ? 1'h0 : _GEN_1849; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1853 = i == 10'h2f3 ? 1'h0 : i == 10'h2f3 | (i == 10'h2f2 | _GEN_1850); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1854 = i == 10'h2f4 ? 1'h0 : _GEN_1853; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1857 = i == 10'h2f5 ? 1'h0 : i == 10'h2f5 | (i == 10'h2f4 | _GEN_1854); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1858 = i == 10'h2f6 ? 1'h0 : _GEN_1857; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1861 = i == 10'h2f7 ? 1'h0 : i == 10'h2f7 | (i == 10'h2f6 | _GEN_1858); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1862 = i == 10'h2f8 ? 1'h0 : _GEN_1861; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1865 = i == 10'h2f9 ? 1'h0 : i == 10'h2f9 | (i == 10'h2f8 | _GEN_1862); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1866 = i == 10'h2fa ? 1'h0 : _GEN_1865; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1869 = i == 10'h2fb ? 1'h0 : i == 10'h2fb | (i == 10'h2fa | _GEN_1866); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1870 = i == 10'h2fc ? 1'h0 : _GEN_1869; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1873 = i == 10'h2fd ? 1'h0 : i == 10'h2fd | (i == 10'h2fc | _GEN_1870); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1874 = i == 10'h2fe ? 1'h0 : _GEN_1873; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1877 = i == 10'h2ff ? 1'h0 : i == 10'h2ff | (i == 10'h2fe | _GEN_1874); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1878 = i == 10'h300 ? 1'h0 : _GEN_1877; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1881 = i == 10'h301 ? 1'h0 : i == 10'h301 | (i == 10'h300 | _GEN_1878); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1882 = i == 10'h302 ? 1'h0 : _GEN_1881; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1885 = i == 10'h303 ? 1'h0 : i == 10'h303 | (i == 10'h302 | _GEN_1882); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1886 = i == 10'h304 ? 1'h0 : _GEN_1885; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1889 = i == 10'h305 ? 1'h0 : i == 10'h305 | (i == 10'h304 | _GEN_1886); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1890 = i == 10'h306 ? 1'h0 : _GEN_1889; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1893 = i == 10'h307 ? 1'h0 : i == 10'h307 | (i == 10'h306 | _GEN_1890); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1894 = i == 10'h308 ? 1'h0 : _GEN_1893; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1897 = i == 10'h309 ? 1'h0 : i == 10'h309 | (i == 10'h308 | _GEN_1894); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1898 = i == 10'h30a ? 1'h0 : _GEN_1897; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1901 = i == 10'h30b ? 1'h0 : i == 10'h30b | (i == 10'h30a | _GEN_1898); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1902 = i == 10'h30c ? 1'h0 : _GEN_1901; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1905 = i == 10'h30d ? 1'h0 : i == 10'h30d | (i == 10'h30c | _GEN_1902); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1906 = i == 10'h30e ? 1'h0 : _GEN_1905; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1909 = i == 10'h30f ? 1'h0 : i == 10'h30f | (i == 10'h30e | _GEN_1906); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1910 = i == 10'h310 ? 1'h0 : _GEN_1909; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1913 = i == 10'h311 ? 1'h0 : i == 10'h311 | (i == 10'h310 | _GEN_1910); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1914 = i == 10'h1 ? 1'h0 : i == 10'h294 | _GEN_1414; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1915 = i == 10'h2 ? 1'h0 : _GEN_1914; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1916 = i == 10'h5 ? 1'h0 : _GEN_1915; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1917 = i == 10'h9 ? 1'h0 : _GEN_1916; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1918 = i == 10'hb ? 1'h0 : _GEN_1917; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1919 = i == 10'h29 ? 1'h0 : _GEN_1918; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1920 = i == 10'h30 ? 1'h0 : _GEN_1919; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1921 = i == 10'h54 ? 1'h0 : _GEN_1920; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1922 = i == 10'h61 ? 1'h0 : _GEN_1921; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1923 = i == 10'haa ? 1'h0 : _GEN_1922; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1924 = i == 10'h156 ? 1'h0 : _GEN_1923; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1925 = i == 10'h188 ? 1'h0 : _GEN_1924; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1926 = i == 10'h2ae ? 1'h0 : _GEN_1925; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1928 = i == 10'h2af ? 1'h0 : i == 10'h2ae | _GEN_1926; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1930 = i == 10'h2b0 ? 1'h0 : i == 10'h2af | _GEN_1928; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1932 = i == 10'h2b1 ? 1'h0 : i == 10'h2b0 | _GEN_1930; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1934 = i == 10'h2b2 ? 1'h0 : i == 10'h2b1 | _GEN_1932; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1936 = i == 10'h2b3 ? 1'h0 : i == 10'h2b2 | _GEN_1934; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1938 = i == 10'h2b4 ? 1'h0 : i == 10'h2b3 | _GEN_1936; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1940 = i == 10'h2b5 ? 1'h0 : i == 10'h2b4 | _GEN_1938; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1942 = i == 10'h2b6 ? 1'h0 : i == 10'h2b5 | _GEN_1940; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1944 = i == 10'h2b7 ? 1'h0 : i == 10'h2b6 | _GEN_1942; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1946 = i == 10'h2b8 ? 1'h0 : i == 10'h2b7 | _GEN_1944; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1948 = i == 10'h2b9 ? 1'h0 : i == 10'h2b8 | _GEN_1946; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1950 = i == 10'h2ba ? 1'h0 : i == 10'h2b9 | _GEN_1948; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1952 = i == 10'h2bb ? 1'h0 : i == 10'h2ba | _GEN_1950; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1954 = i == 10'h2bc ? 1'h0 : i == 10'h2bb | _GEN_1952; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1956 = i == 10'h2bd ? 1'h0 : i == 10'h2bc | _GEN_1954; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1958 = i == 10'h2be ? 1'h0 : i == 10'h2bd | _GEN_1956; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1960 = i == 10'h2bf ? 1'h0 : i == 10'h2be | _GEN_1958; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1962 = i == 10'h2c0 ? 1'h0 : i == 10'h2bf | _GEN_1960; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1964 = i == 10'h2c1 ? 1'h0 : i == 10'h2c0 | _GEN_1962; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1966 = i == 10'h2c2 ? 1'h0 : i == 10'h2c1 | _GEN_1964; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1968 = i == 10'h2c3 ? 1'h0 : i == 10'h2c2 | _GEN_1966; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1970 = i == 10'h2c4 ? 1'h0 : i == 10'h2c3 | _GEN_1968; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1972 = i == 10'h2c5 ? 1'h0 : i == 10'h2c4 | _GEN_1970; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1974 = i == 10'h2c6 ? 1'h0 : i == 10'h2c5 | _GEN_1972; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1976 = i == 10'h2c7 ? 1'h0 : i == 10'h2c6 | _GEN_1974; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1978 = i == 10'h2c8 ? 1'h0 : i == 10'h2c7 | _GEN_1976; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1980 = i == 10'h2c9 ? 1'h0 : i == 10'h2c8 | _GEN_1978; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1982 = i == 10'h2ca ? 1'h0 : i == 10'h2c9 | _GEN_1980; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1984 = i == 10'h2cb ? 1'h0 : i == 10'h2ca | _GEN_1982; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1986 = i == 10'h2cc ? 1'h0 : i == 10'h2cb | _GEN_1984; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1988 = i == 10'h2cd ? 1'h0 : i == 10'h2cc | _GEN_1986; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1990 = i == 10'h2ce ? 1'h0 : i == 10'h2cd | _GEN_1988; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1992 = i == 10'h2cf ? 1'h0 : i == 10'h2ce | _GEN_1990; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1994 = i == 10'h2d0 ? 1'h0 : i == 10'h2cf | _GEN_1992; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1996 = i == 10'h2d1 ? 1'h0 : i == 10'h2d0 | _GEN_1994; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1998 = i == 10'h2d2 ? 1'h0 : i == 10'h2d1 | _GEN_1996; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2000 = i == 10'h2d3 ? 1'h0 : i == 10'h2d2 | _GEN_1998; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2002 = i == 10'h2d4 ? 1'h0 : i == 10'h2d3 | _GEN_2000; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2004 = i == 10'h2d5 ? 1'h0 : i == 10'h2d4 | _GEN_2002; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2006 = i == 10'h2d6 ? 1'h0 : i == 10'h2d5 | _GEN_2004; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2008 = i == 10'h2d7 ? 1'h0 : i == 10'h2d6 | _GEN_2006; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2010 = i == 10'h2d8 ? 1'h0 : i == 10'h2d7 | _GEN_2008; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2012 = i == 10'h2d9 ? 1'h0 : i == 10'h2d8 | _GEN_2010; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2014 = i == 10'h2da ? 1'h0 : i == 10'h2d9 | _GEN_2012; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2016 = i == 10'h2db ? 1'h0 : i == 10'h2da | _GEN_2014; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2018 = i == 10'h2dc ? 1'h0 : i == 10'h2db | _GEN_2016; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2020 = i == 10'h2dd ? 1'h0 : i == 10'h2dc | _GEN_2018; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2022 = i == 10'h2de ? 1'h0 : i == 10'h2dd | _GEN_2020; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2024 = i == 10'h2df ? 1'h0 : i == 10'h2de | _GEN_2022; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2026 = i == 10'h2e0 ? 1'h0 : i == 10'h2df | _GEN_2024; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2028 = i == 10'h2e1 ? 1'h0 : i == 10'h2e0 | _GEN_2026; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2030 = i == 10'h2e2 ? 1'h0 : i == 10'h2e1 | _GEN_2028; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2032 = i == 10'h2e3 ? 1'h0 : i == 10'h2e2 | _GEN_2030; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2034 = i == 10'h2e4 ? 1'h0 : i == 10'h2e3 | _GEN_2032; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2036 = i == 10'h2e5 ? 1'h0 : i == 10'h2e4 | _GEN_2034; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2038 = i == 10'h2e6 ? 1'h0 : i == 10'h2e5 | _GEN_2036; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2040 = i == 10'h2e7 ? 1'h0 : i == 10'h2e6 | _GEN_2038; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2042 = i == 10'h2e8 ? 1'h0 : i == 10'h2e7 | _GEN_2040; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2044 = i == 10'h2e9 ? 1'h0 : i == 10'h2e8 | _GEN_2042; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2046 = i == 10'h2ea ? 1'h0 : i == 10'h2e9 | _GEN_2044; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2048 = i == 10'h2eb ? 1'h0 : i == 10'h2ea | _GEN_2046; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2050 = i == 10'h2ec ? 1'h0 : i == 10'h2eb | _GEN_2048; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2052 = i == 10'h2ed ? 1'h0 : i == 10'h2ec | _GEN_2050; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2054 = i == 10'h2ee ? 1'h0 : i == 10'h2ed | _GEN_2052; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2056 = i == 10'h2ef ? 1'h0 : i == 10'h2ee | _GEN_2054; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2058 = i == 10'h2f0 ? 1'h0 : i == 10'h2ef | _GEN_2056; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2060 = i == 10'h2f1 ? 1'h0 : i == 10'h2f0 | _GEN_2058; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2062 = i == 10'h2f2 ? 1'h0 : i == 10'h2f1 | _GEN_2060; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2064 = i == 10'h2f3 ? 1'h0 : i == 10'h2f2 | _GEN_2062; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2066 = i == 10'h2f4 ? 1'h0 : i == 10'h2f3 | _GEN_2064; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2068 = i == 10'h2f5 ? 1'h0 : i == 10'h2f4 | _GEN_2066; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2070 = i == 10'h2f6 ? 1'h0 : i == 10'h2f5 | _GEN_2068; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2072 = i == 10'h2f7 ? 1'h0 : i == 10'h2f6 | _GEN_2070; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2074 = i == 10'h2f8 ? 1'h0 : i == 10'h2f7 | _GEN_2072; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2076 = i == 10'h2f9 ? 1'h0 : i == 10'h2f8 | _GEN_2074; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2078 = i == 10'h2fa ? 1'h0 : i == 10'h2f9 | _GEN_2076; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2080 = i == 10'h2fb ? 1'h0 : i == 10'h2fa | _GEN_2078; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2082 = i == 10'h2fc ? 1'h0 : i == 10'h2fb | _GEN_2080; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2084 = i == 10'h2fd ? 1'h0 : i == 10'h2fc | _GEN_2082; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2086 = i == 10'h2fe ? 1'h0 : i == 10'h2fd | _GEN_2084; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2088 = i == 10'h2ff ? 1'h0 : i == 10'h2fe | _GEN_2086; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2090 = i == 10'h300 ? 1'h0 : i == 10'h2ff | _GEN_2088; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2092 = i == 10'h301 ? 1'h0 : i == 10'h300 | _GEN_2090; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2094 = i == 10'h302 ? 1'h0 : i == 10'h301 | _GEN_2092; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2096 = i == 10'h303 ? 1'h0 : i == 10'h302 | _GEN_2094; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2098 = i == 10'h304 ? 1'h0 : i == 10'h303 | _GEN_2096; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2100 = i == 10'h305 ? 1'h0 : i == 10'h304 | _GEN_2098; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2102 = i == 10'h306 ? 1'h0 : i == 10'h305 | _GEN_2100; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2104 = i == 10'h307 ? 1'h0 : i == 10'h306 | _GEN_2102; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2106 = i == 10'h308 ? 1'h0 : i == 10'h307 | _GEN_2104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2108 = i == 10'h309 ? 1'h0 : i == 10'h308 | _GEN_2106; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2110 = i == 10'h30a ? 1'h0 : i == 10'h309 | _GEN_2108; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2112 = i == 10'h30b ? 1'h0 : i == 10'h30a | _GEN_2110; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2114 = i == 10'h30c ? 1'h0 : i == 10'h30b | _GEN_2112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2116 = i == 10'h30d ? 1'h0 : i == 10'h30c | _GEN_2114; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2118 = i == 10'h30e ? 1'h0 : i == 10'h30d | _GEN_2116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2120 = i == 10'h30f ? 1'h0 : i == 10'h30e | _GEN_2118; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2122 = i == 10'h310 ? 1'h0 : i == 10'h30f | _GEN_2120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2124 = i == 10'h311 ? 1'h0 : i == 10'h310 | _GEN_2122; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2126 = i == 10'h0 ? 1'h0 : _GEN_1431; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2130 = i == 10'h17 ? 1'h0 : i == 10'hb | (i == 10'h5 | (i == 10'h2 | _GEN_2126)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2131 = i == 10'h30 ? 1'h0 : _GEN_2130; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2133 = i == 10'hc5 ? 1'h0 : i == 10'h62 | _GEN_2131; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2134 = i == 10'hc5 | _GEN_2133; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2135 = i == 10'h0 ? 1'h0 : _GEN_1471; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2139 = i == 10'h2f ? 1'h0 : i == 10'h18 | (i == 10'h5 | (i == 10'h2 | _GEN_2135)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2141 = i == 10'h31 ? 1'h0 : i == 10'h30 | _GEN_2139; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2143 = i == 10'h62 ? 1'h0 : i == 10'h60 | _GEN_2141; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2145 = i == 10'hc1 ? 1'h0 : i == 10'h64 | _GEN_2143; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2148 = i == 10'hc5 ? 1'h0 : i == 10'hc5 | (i == 10'hc1 | _GEN_2145); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2149 = i == 10'hc9 ? 1'h0 : _GEN_2148; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2150 = i == 10'hc9 | _GEN_2149; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2151 = i == 10'h0 ? 1'h0 : _GEN_1532; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2152 = i == 10'h2 ? 1'h0 : _GEN_2151; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2153 = i == 10'h5 ? 1'h0 : _GEN_2152; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2154 = i == 10'h18 ? 1'h0 : _GEN_2153; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2156 = i == 10'h60 ? 1'h0 : i == 10'h5f | _GEN_2154; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2158 = i == 10'h62 ? 1'h0 : i == 10'h61 | _GEN_2156; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2160 = i == 10'h64 ? 1'h0 : i == 10'h63 | _GEN_2158; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2161 = i == 10'hbf ? 1'h0 : _GEN_2160; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2164 = i == 10'hc1 ? 1'h0 : i == 10'hc1 | (i == 10'hbf | _GEN_2161); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2165 = i == 10'hc3 ? 1'h0 : _GEN_2164; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2168 = i == 10'hc5 ? 1'h0 : i == 10'hc5 | (i == 10'hc3 | _GEN_2165); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2169 = i == 10'hc7 ? 1'h0 : _GEN_2168; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2173 = i == 10'h1 ? 1'h0 : _GEN_1623; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2174 = i == 10'h2 ? 1'h0 : _GEN_2173; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2175 = i == 10'h4 ? 1'h0 : _GEN_2174; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2176 = i == 10'h5 ? 1'h0 : _GEN_2175; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2177 = i == 10'ha ? 1'h0 : _GEN_2176; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2178 = i == 10'h16 ? 1'h0 : _GEN_2177; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2179 = i == 10'h18 ? 1'h0 : _GEN_2178; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2180 = i == 10'h2e ? 1'h0 : _GEN_2179; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2181 = i == 10'h5e ? 1'h0 : _GEN_2180; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2182 = i == 10'h64 ? 1'h0 : _GEN_2181; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2183 = i == 10'hbe ? 1'h0 : _GEN_2182; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2186 = i == 10'hbf ? 1'h0 : i == 10'hbf | (i == 10'hbe | _GEN_2183); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2187 = i == 10'hc0 ? 1'h0 : _GEN_2186; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2190 = i == 10'hc1 ? 1'h0 : i == 10'hc1 | (i == 10'hc0 | _GEN_2187); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2191 = i == 10'hc2 ? 1'h0 : _GEN_2190; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2194 = i == 10'hc3 ? 1'h0 : i == 10'hc3 | (i == 10'hc2 | _GEN_2191); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2195 = i == 10'hc4 ? 1'h0 : _GEN_2194; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2198 = i == 10'hc5 ? 1'h0 : i == 10'hc5 | (i == 10'hc4 | _GEN_2195); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2199 = i == 10'hc6 ? 1'h0 : _GEN_2198; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2202 = i == 10'hc7 ? 1'h0 : i == 10'hc7 | (i == 10'hc6 | _GEN_2199); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2203 = i == 10'hc8 ? 1'h0 : _GEN_2202; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2207 = i == 10'h1 ? 1'h0 : _GEN_1755; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2209 = i == 10'h4 ? 1'h0 : i == 10'h2 | _GEN_2207; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2211 = i == 10'ha ? 1'h0 : i == 10'h5 | _GEN_2209; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2212 = i == 10'h16 ? 1'h0 : _GEN_2211; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2214 = i == 10'h2e ? 1'h0 : i == 10'h18 | _GEN_2212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2215 = i == 10'h5e ? 1'h0 : _GEN_2214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2218 = i == 10'hbe ? 1'h0 : i == 10'hbe | (i == 10'h64 | _GEN_2215); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2220 = i == 10'hbf ? 1'h0 : i == 10'hbf | _GEN_2218; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2222 = i == 10'hc0 ? 1'h0 : i == 10'hc0 | _GEN_2220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2224 = i == 10'hc1 ? 1'h0 : i == 10'hc1 | _GEN_2222; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2226 = i == 10'hc2 ? 1'h0 : i == 10'hc2 | _GEN_2224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2228 = i == 10'hc3 ? 1'h0 : i == 10'hc3 | _GEN_2226; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2230 = i == 10'hc4 ? 1'h0 : i == 10'hc4 | _GEN_2228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2232 = i == 10'hc5 ? 1'h0 : i == 10'hc5 | _GEN_2230; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2234 = i == 10'hc6 ? 1'h0 : i == 10'hc6 | _GEN_2232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2236 = i == 10'hc7 ? 1'h0 : i == 10'hc7 | _GEN_2234; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2238 = i == 10'hc8 ? 1'h0 : i == 10'hc8 | _GEN_2236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2241 = i == 10'h1 ? 1'h0 : _GEN_1913; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2242 = i == 10'h2 ? 1'h0 : _GEN_2241; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2243 = i == 10'h4 ? 1'h0 : _GEN_2242; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2244 = i == 10'h5 ? 1'h0 : _GEN_2243; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2245 = i == 10'ha ? 1'h0 : _GEN_2244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2246 = i == 10'h16 ? 1'h0 : _GEN_2245; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2247 = i == 10'h18 ? 1'h0 : _GEN_2246; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2248 = i == 10'h2e ? 1'h0 : _GEN_2247; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2249 = i == 10'h64 ? 1'h0 : _GEN_2248; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2250 = i == 10'hbd ? 1'h0 : _GEN_2249; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2251 = i == 10'h17c ? 1'h0 : _GEN_2250; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2253 = i == 10'h17d ? 1'h0 : i == 10'h17c | _GEN_2251; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2255 = i == 10'h17e ? 1'h0 : i == 10'h17d | _GEN_2253; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2257 = i == 10'h17f ? 1'h0 : i == 10'h17e | _GEN_2255; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2259 = i == 10'h180 ? 1'h0 : i == 10'h17f | _GEN_2257; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2261 = i == 10'h181 ? 1'h0 : i == 10'h180 | _GEN_2259; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2263 = i == 10'h182 ? 1'h0 : i == 10'h181 | _GEN_2261; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2265 = i == 10'h183 ? 1'h0 : i == 10'h182 | _GEN_2263; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2267 = i == 10'h184 ? 1'h0 : i == 10'h183 | _GEN_2265; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2269 = i == 10'h185 ? 1'h0 : i == 10'h184 | _GEN_2267; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2271 = i == 10'h186 ? 1'h0 : i == 10'h185 | _GEN_2269; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2273 = i == 10'h187 ? 1'h0 : i == 10'h186 | _GEN_2271; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2275 = i == 10'h188 ? 1'h0 : i == 10'h187 | _GEN_2273; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2277 = i == 10'h189 ? 1'h0 : i == 10'h188 | _GEN_2275; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2279 = i == 10'h18a ? 1'h0 : i == 10'h189 | _GEN_2277; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2281 = i == 10'h18b ? 1'h0 : i == 10'h18a | _GEN_2279; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2283 = i == 10'h18c ? 1'h0 : i == 10'h18b | _GEN_2281; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2285 = i == 10'h18d ? 1'h0 : i == 10'h18c | _GEN_2283; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2287 = i == 10'h18e ? 1'h0 : i == 10'h18d | _GEN_2285; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2289 = i == 10'h18f ? 1'h0 : i == 10'h18e | _GEN_2287; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2291 = i == 10'h190 ? 1'h0 : i == 10'h18f | _GEN_2289; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2293 = i == 10'h191 ? 1'h0 : i == 10'h190 | _GEN_2291; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2295 = i == 10'h192 ? 1'h0 : i == 10'h191 | _GEN_2293; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2297 = i == 10'h193 ? 1'h0 : i == 10'h192 | _GEN_2295; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2299 = i == 10'h194 ? 1'h0 : i == 10'h193 | _GEN_2297; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2300 = i == 10'h194 | _GEN_2299; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2301 = i == 10'h1 ? 1'h0 : i == 10'h311 | _GEN_2124; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2302 = i == 10'h2 ? 1'h0 : _GEN_2301; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2303 = i == 10'h4 ? 1'h0 : _GEN_2302; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2304 = i == 10'h5 ? 1'h0 : _GEN_2303; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2305 = i == 10'ha ? 1'h0 : _GEN_2304; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2306 = i == 10'h16 ? 1'h0 : _GEN_2305; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2307 = i == 10'h18 ? 1'h0 : _GEN_2306; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2308 = i == 10'h2e ? 1'h0 : _GEN_2307; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2309 = i == 10'h64 ? 1'h0 : _GEN_2308; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2310 = i == 10'hbd ? 1'h0 : _GEN_2309; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2311 = i == 10'h2f9 ? 1'h0 : _GEN_2310; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2313 = i == 10'h2fa ? 1'h0 : i == 10'h2f9 | _GEN_2311; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2315 = i == 10'h2fb ? 1'h0 : i == 10'h2fa | _GEN_2313; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2317 = i == 10'h2fc ? 1'h0 : i == 10'h2fb | _GEN_2315; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2319 = i == 10'h2fd ? 1'h0 : i == 10'h2fc | _GEN_2317; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2321 = i == 10'h2fe ? 1'h0 : i == 10'h2fd | _GEN_2319; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2323 = i == 10'h2ff ? 1'h0 : i == 10'h2fe | _GEN_2321; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2325 = i == 10'h300 ? 1'h0 : i == 10'h2ff | _GEN_2323; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2327 = i == 10'h301 ? 1'h0 : i == 10'h300 | _GEN_2325; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2329 = i == 10'h302 ? 1'h0 : i == 10'h301 | _GEN_2327; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2331 = i == 10'h303 ? 1'h0 : i == 10'h302 | _GEN_2329; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2333 = i == 10'h304 ? 1'h0 : i == 10'h303 | _GEN_2331; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2335 = i == 10'h305 ? 1'h0 : i == 10'h304 | _GEN_2333; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2337 = i == 10'h306 ? 1'h0 : i == 10'h305 | _GEN_2335; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2339 = i == 10'h307 ? 1'h0 : i == 10'h306 | _GEN_2337; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2341 = i == 10'h308 ? 1'h0 : i == 10'h307 | _GEN_2339; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2343 = i == 10'h309 ? 1'h0 : i == 10'h308 | _GEN_2341; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2345 = i == 10'h30a ? 1'h0 : i == 10'h309 | _GEN_2343; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2347 = i == 10'h30b ? 1'h0 : i == 10'h30a | _GEN_2345; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2349 = i == 10'h30c ? 1'h0 : i == 10'h30b | _GEN_2347; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2351 = i == 10'h30d ? 1'h0 : i == 10'h30c | _GEN_2349; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2353 = i == 10'h30e ? 1'h0 : i == 10'h30d | _GEN_2351; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2355 = i == 10'h30f ? 1'h0 : i == 10'h30e | _GEN_2353; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2357 = i == 10'h310 ? 1'h0 : i == 10'h30f | _GEN_2355; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2359 = i == 10'h311 ? 1'h0 : i == 10'h310 | _GEN_2357; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2361 = i == 10'h312 ? 1'h0 : i == 10'h311 | _GEN_2359; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2363 = i == 10'h313 ? 1'h0 : i == 10'h312 | _GEN_2361; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2365 = i == 10'h314 ? 1'h0 : i == 10'h313 | _GEN_2363; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2367 = i == 10'h315 ? 1'h0 : i == 10'h314 | _GEN_2365; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2369 = i == 10'h316 ? 1'h0 : i == 10'h315 | _GEN_2367; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2371 = i == 10'h317 ? 1'h0 : i == 10'h316 | _GEN_2369; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2373 = i == 10'h318 ? 1'h0 : i == 10'h317 | _GEN_2371; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2375 = i == 10'h319 ? 1'h0 : i == 10'h318 | _GEN_2373; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2377 = i == 10'h31a ? 1'h0 : i == 10'h319 | _GEN_2375; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2379 = i == 10'h31b ? 1'h0 : i == 10'h31a | _GEN_2377; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2381 = i == 10'h31c ? 1'h0 : i == 10'h31b | _GEN_2379; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2383 = i == 10'h31d ? 1'h0 : i == 10'h31c | _GEN_2381; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2385 = i == 10'h31e ? 1'h0 : i == 10'h31d | _GEN_2383; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2387 = i == 10'h31f ? 1'h0 : i == 10'h31e | _GEN_2385; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2389 = i == 10'h320 ? 1'h0 : i == 10'h31f | _GEN_2387; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2391 = i == 10'h321 ? 1'h0 : i == 10'h320 | _GEN_2389; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2393 = i == 10'h322 ? 1'h0 : i == 10'h321 | _GEN_2391; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2395 = i == 10'h323 ? 1'h0 : i == 10'h322 | _GEN_2393; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2397 = i == 10'h324 ? 1'h0 : i == 10'h323 | _GEN_2395; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2399 = i == 10'h325 ? 1'h0 : i == 10'h324 | _GEN_2397; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2401 = i == 10'h326 ? 1'h0 : i == 10'h325 | _GEN_2399; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2403 = i == 10'h327 ? 1'h0 : i == 10'h326 | _GEN_2401; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2405 = i == 10'h328 ? 1'h0 : i == 10'h327 | _GEN_2403; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2407 = i == 10'h329 ? 1'h0 : i == 10'h328 | _GEN_2405; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2409 = i == 10'h32a ? 1'h0 : i == 10'h329 | _GEN_2407; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2410 = i == 10'h32a | _GEN_2409; // @[lut_mem_online.scala 235:34 239:30]
  wire  _T_2414 = counter < 5'h11; // @[lut_mem_online.scala 250:22]
  wire  _T_2416 = counter >= 5'ha; // @[lut_mem_online.scala 258:30]
  wire [4:0] _outResult_T_1 = counter - 5'ha; // @[lut_mem_online.scala 260:41]
  wire  _GEN_2419 = 4'h1 == _outResult_T_1[3:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2420 = 4'h2 == _outResult_T_1[3:0] ? buffer_2 : _GEN_2419; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2421 = 4'h3 == _outResult_T_1[3:0] ? buffer_3 : _GEN_2420; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2422 = 4'h4 == _outResult_T_1[3:0] ? buffer_4 : _GEN_2421; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2423 = 4'h5 == _outResult_T_1[3:0] ? buffer_5 : _GEN_2422; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2424 = 4'h6 == _outResult_T_1[3:0] ? buffer_6 : _GEN_2423; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2425 = 4'h7 == _outResult_T_1[3:0] ? 1'h0 : _GEN_2424; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2426 = 4'h8 == _outResult_T_1[3:0] ? 1'h0 : _GEN_2425; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_2427 = 4'h9 == _outResult_T_1[3:0] ? 1'h0 : _GEN_2426; // @[lut_mem_online.scala 260:{23,23}]
  wire  _T_2420 = ~reset; // @[lut_mem_online.scala 263:21]
  wire  _GEN_2429 = counter >= 5'ha ? _GEN_2427 : outResult; // @[lut_mem_online.scala 258:42 260:23 215:26]
  wire  _GEN_2431 = _T_2 ? 1'h0 : _GEN_2429; // @[lut_mem_online.scala 255:35 257:23]
  wire  _T_2421 = i < 10'h1ff; // @[lut_mem_online.scala 274:18]
  wire [11:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 284:24]
  wire [11:0] _i_T_2 = _i_T + 12'h1; // @[lut_mem_online.scala 284:28]
  wire [11:0] _i_T_5 = _i_T + 12'h2; // @[lut_mem_online.scala 286:28]
  wire [11:0] _GEN_2432 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 285:45 286:17 206:18]
  wire [11:0] _GEN_2433 = ~io_inputBit ? _i_T_2 : _GEN_2432; // @[lut_mem_online.scala 283:39 284:17]
  wire  _T_2426 = i < 10'h3ff; // @[lut_mem_online.scala 289:24]
  wire [9:0] _GEN_2434 = i < 10'h3ff ? 10'h3ff : i; // @[lut_mem_online.scala 289:63 297:15 206:18]
  wire [11:0] _GEN_2435 = i < 10'h1ff ? _GEN_2433 : {{2'd0}, _GEN_2434}; // @[lut_mem_online.scala 274:61]
  wire [4:0] _counter_T_1 = counter + 5'h1; // @[lut_mem_online.scala 300:30]
  wire  _GEN_2437 = counter < 5'h11 & _GEN_2431; // @[lut_mem_online.scala 250:52 304:21]
  wire [11:0] _GEN_2438 = counter < 5'h11 ? _GEN_2435 : {{2'd0}, i}; // @[lut_mem_online.scala 206:18 250:52]
  wire  _GEN_2461 = io_start & _GEN_2437; // @[lut_mem_online.scala 220:29 327:15]
  wire [11:0] _GEN_2462 = io_start ? _GEN_2438 : 12'h0; // @[lut_mem_online.scala 220:29 325:7]
  wire [11:0] _GEN_2465 = reset ? 12'h0 : _GEN_2462; // @[lut_mem_online.scala 206:{18,18}]
  wire  _GEN_2466 = io_start & _T_2414; // @[lut_mem_online.scala 263:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 334:16]
  always @(posedge clock) begin
    i <= _GEN_2465[9:0]; // @[lut_mem_online.scala 206:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        buffer_0 <= _GEN_2134;
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        buffer_1 <= _GEN_2150;
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 235:34]
          buffer_2 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_2 <= i == 10'hc9 | (i == 10'hc7 | _GEN_2169);
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 235:34]
          buffer_3 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_3 <= i == 10'hc9 | (i == 10'hc8 | _GEN_2203);
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 235:34]
          buffer_4 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_4 <= i == 10'hc9 | _GEN_2238;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        buffer_5 <= _GEN_2300;
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 232:36]
        buffer_6 <= _GEN_2410;
      end
    end
    if (reset) begin // @[lut_mem_online.scala 212:24]
      counter <= 5'h0; // @[lut_mem_online.scala 212:24]
    end else if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h11) begin // @[lut_mem_online.scala 250:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 300:19]
      end
    end else begin
      counter <= 5'h0; // @[lut_mem_online.scala 326:13]
    end
    if (reset) begin // @[lut_mem_online.scala 215:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 215:26]
    end else begin
      outResult <= _GEN_2461;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_2414 & ~_T_2 & _T_2416 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 263:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2466 & _T_2421 & _T_2420) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 277:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2466 & ~_T_2421 & _T_2426 & _T_2420) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 292:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
