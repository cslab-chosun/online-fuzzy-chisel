module LutMembershipFunctionOnline_9(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [9:0] i; // @[lut_mem_online.scala 205:18]
  reg  buffer_0; // @[lut_mem_online.scala 209:19]
  reg  buffer_1; // @[lut_mem_online.scala 209:19]
  reg  buffer_2; // @[lut_mem_online.scala 209:19]
  reg  buffer_3; // @[lut_mem_online.scala 209:19]
  reg  buffer_4; // @[lut_mem_online.scala 209:19]
  reg  buffer_5; // @[lut_mem_online.scala 209:19]
  reg  buffer_6; // @[lut_mem_online.scala 209:19]
  reg [4:0] counter; // @[lut_mem_online.scala 211:24]
  reg  outResult; // @[lut_mem_online.scala 214:26]
  wire  _T_2 = counter < 5'ha; // @[lut_mem_online.scala 231:22]
  wire  _GEN_0 = io_inputBit ? 1'h0 : buffer_0; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_1 = i == 10'h0 ? _GEN_0 : buffer_0; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_2 = io_inputBit ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3 = i == 10'h1 ? _GEN_2 : _GEN_1; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4 = io_inputBit ? 1'h0 : _GEN_3; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5 = i == 10'h3 ? _GEN_4 : _GEN_3; // @[lut_mem_online.scala 234:34]
  wire  _T_10 = ~io_inputBit; // @[lut_mem_online.scala 236:32]
  wire  _GEN_6 = ~io_inputBit | _GEN_5; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_7 = i == 10'h7 ? _GEN_6 : _GEN_5; // @[lut_mem_online.scala 234:34]
  wire  _GEN_8 = ~io_inputBit | _GEN_7; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_9 = i == 10'h10 ? _GEN_8 : _GEN_7; // @[lut_mem_online.scala 234:34]
  wire  _GEN_10 = ~io_inputBit | _GEN_9; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_11 = i == 10'h22 ? _GEN_10 : _GEN_9; // @[lut_mem_online.scala 234:34]
  wire  _GEN_12 = io_inputBit ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_13 = i == 10'h22 ? _GEN_12 : _GEN_11; // @[lut_mem_online.scala 234:34]
  wire  _GEN_14 = io_inputBit ? 1'h0 : buffer_1; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_15 = i == 10'h0 ? _GEN_14 : buffer_1; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_16 = io_inputBit ? 1'h0 : _GEN_15; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_17 = i == 10'h1 ? _GEN_16 : _GEN_15; // @[lut_mem_online.scala 234:34]
  wire  _GEN_18 = ~io_inputBit | _GEN_17; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_19 = i == 10'h7 ? _GEN_18 : _GEN_17; // @[lut_mem_online.scala 234:34]
  wire  _GEN_20 = io_inputBit ? 1'h0 : _GEN_19; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_21 = i == 10'h8 ? _GEN_20 : _GEN_19; // @[lut_mem_online.scala 234:34]
  wire  _GEN_22 = io_inputBit ? 1'h0 : _GEN_21; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_23 = i == 10'h11 ? _GEN_22 : _GEN_21; // @[lut_mem_online.scala 234:34]
  wire  _GEN_24 = ~io_inputBit | _GEN_23; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_25 = i == 10'h21 ? _GEN_24 : _GEN_23; // @[lut_mem_online.scala 234:34]
  wire  _GEN_26 = ~io_inputBit ? 1'h0 : _GEN_25; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_27 = i == 10'h22 ? _GEN_26 : _GEN_25; // @[lut_mem_online.scala 234:34]
  wire  _GEN_28 = io_inputBit | _GEN_27; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_29 = i == 10'h22 ? _GEN_28 : _GEN_27; // @[lut_mem_online.scala 234:34]
  wire  _GEN_30 = io_inputBit ? 1'h0 : _GEN_29; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_31 = i == 10'h23 ? _GEN_30 : _GEN_29; // @[lut_mem_online.scala 234:34]
  wire  _GEN_32 = io_inputBit ? 1'h0 : _GEN_31; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_33 = i == 10'h44 ? _GEN_32 : _GEN_31; // @[lut_mem_online.scala 234:34]
  wire  _GEN_34 = ~io_inputBit | _GEN_33; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_35 = i == 10'h47 ? _GEN_34 : _GEN_33; // @[lut_mem_online.scala 234:34]
  wire  _GEN_36 = io_inputBit ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_37 = i == 10'h47 ? _GEN_36 : _GEN_35; // @[lut_mem_online.scala 234:34]
  wire  _GEN_38 = ~io_inputBit | _GEN_37; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_39 = i == 10'h89 ? _GEN_38 : _GEN_37; // @[lut_mem_online.scala 234:34]
  wire  _GEN_40 = io_inputBit ? 1'h0 : _GEN_39; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_41 = i == 10'h89 ? _GEN_40 : _GEN_39; // @[lut_mem_online.scala 234:34]
  wire  _GEN_42 = io_inputBit ? 1'h0 : buffer_2; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_43 = i == 10'h0 ? _GEN_42 : buffer_2; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_44 = io_inputBit ? 1'h0 : _GEN_43; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_45 = i == 10'h1 ? _GEN_44 : _GEN_43; // @[lut_mem_online.scala 234:34]
  wire  _GEN_46 = ~io_inputBit ? 1'h0 : _GEN_45; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_47 = i == 10'h7 ? _GEN_46 : _GEN_45; // @[lut_mem_online.scala 234:34]
  wire  _GEN_48 = io_inputBit ? 1'h0 : _GEN_47; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_49 = i == 10'h8 ? _GEN_48 : _GEN_47; // @[lut_mem_online.scala 234:34]
  wire  _GEN_50 = io_inputBit ? 1'h0 : _GEN_49; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_51 = i == 10'h11 ? _GEN_50 : _GEN_49; // @[lut_mem_online.scala 234:34]
  wire  _GEN_52 = ~io_inputBit ? 1'h0 : _GEN_51; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_53 = i == 10'h21 ? _GEN_52 : _GEN_51; // @[lut_mem_online.scala 234:34]
  wire  _GEN_54 = io_inputBit | _GEN_53; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_55 = i == 10'h44 ? _GEN_54 : _GEN_53; // @[lut_mem_online.scala 234:34]
  wire  _GEN_56 = io_inputBit ? 1'h0 : _GEN_55; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_57 = i == 10'h45 ? _GEN_56 : _GEN_55; // @[lut_mem_online.scala 234:34]
  wire  _GEN_58 = ~io_inputBit | _GEN_57; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_59 = i == 10'h46 ? _GEN_58 : _GEN_57; // @[lut_mem_online.scala 234:34]
  wire  _GEN_60 = ~io_inputBit ? 1'h0 : _GEN_59; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_61 = i == 10'h47 ? _GEN_60 : _GEN_59; // @[lut_mem_online.scala 234:34]
  wire  _GEN_62 = io_inputBit | _GEN_61; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_63 = i == 10'h47 ? _GEN_62 : _GEN_61; // @[lut_mem_online.scala 234:34]
  wire  _GEN_64 = io_inputBit ? 1'h0 : _GEN_63; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_65 = i == 10'h48 ? _GEN_64 : _GEN_63; // @[lut_mem_online.scala 234:34]
  wire  _GEN_66 = ~io_inputBit ? 1'h0 : _GEN_65; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_67 = i == 10'h89 ? _GEN_66 : _GEN_65; // @[lut_mem_online.scala 234:34]
  wire  _GEN_68 = io_inputBit | _GEN_67; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_69 = i == 10'h89 ? _GEN_68 : _GEN_67; // @[lut_mem_online.scala 234:34]
  wire  _GEN_70 = ~io_inputBit | _GEN_69; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_71 = i == 10'h8b ? _GEN_70 : _GEN_69; // @[lut_mem_online.scala 234:34]
  wire  _GEN_72 = io_inputBit ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_73 = i == 10'h8b ? _GEN_72 : _GEN_71; // @[lut_mem_online.scala 234:34]
  wire  _GEN_74 = ~io_inputBit | _GEN_73; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_75 = i == 10'h8e ? _GEN_74 : _GEN_73; // @[lut_mem_online.scala 234:34]
  wire  _GEN_76 = io_inputBit ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_77 = i == 10'h8e ? _GEN_76 : _GEN_75; // @[lut_mem_online.scala 234:34]
  wire  _GEN_78 = ~io_inputBit | _GEN_77; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_79 = i == 10'h91 ? _GEN_78 : _GEN_77; // @[lut_mem_online.scala 234:34]
  wire  _GEN_80 = io_inputBit ? 1'h0 : _GEN_79; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_81 = i == 10'h91 ? _GEN_80 : _GEN_79; // @[lut_mem_online.scala 234:34]
  wire  _GEN_82 = io_inputBit ? 1'h0 : buffer_3; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_83 = i == 10'h0 ? _GEN_82 : buffer_3; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_84 = io_inputBit ? 1'h0 : _GEN_83; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_85 = i == 10'h1 ? _GEN_84 : _GEN_83; // @[lut_mem_online.scala 234:34]
  wire  _GEN_86 = ~io_inputBit ? 1'h0 : _GEN_85; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_87 = i == 10'h7 ? _GEN_86 : _GEN_85; // @[lut_mem_online.scala 234:34]
  wire  _GEN_88 = io_inputBit ? 1'h0 : _GEN_87; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_89 = i == 10'h8 ? _GEN_88 : _GEN_87; // @[lut_mem_online.scala 234:34]
  wire  _GEN_90 = io_inputBit ? 1'h0 : _GEN_89; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_91 = i == 10'h11 ? _GEN_90 : _GEN_89; // @[lut_mem_online.scala 234:34]
  wire  _GEN_92 = ~io_inputBit ? 1'h0 : _GEN_91; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_93 = i == 10'h21 ? _GEN_92 : _GEN_91; // @[lut_mem_online.scala 234:34]
  wire  _GEN_94 = io_inputBit ? 1'h0 : _GEN_93; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_95 = i == 10'h45 ? _GEN_94 : _GEN_93; // @[lut_mem_online.scala 234:34]
  wire  _GEN_96 = io_inputBit | _GEN_95; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_97 = i == 10'h47 ? _GEN_96 : _GEN_95; // @[lut_mem_online.scala 234:34]
  wire  _GEN_98 = ~io_inputBit ? 1'h0 : _GEN_97; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_99 = i == 10'h89 ? _GEN_98 : _GEN_97; // @[lut_mem_online.scala 234:34]
  wire  _GEN_100 = io_inputBit | _GEN_99; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_101 = i == 10'h89 ? _GEN_100 : _GEN_99; // @[lut_mem_online.scala 234:34]
  wire  _GEN_102 = ~io_inputBit | _GEN_101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_103 = i == 10'h8a ? _GEN_102 : _GEN_101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_104 = io_inputBit ? 1'h0 : _GEN_103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_105 = i == 10'h8a ? _GEN_104 : _GEN_103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_106 = ~io_inputBit ? 1'h0 : _GEN_105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_107 = i == 10'h8b ? _GEN_106 : _GEN_105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_108 = io_inputBit | _GEN_107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_109 = i == 10'h8b ? _GEN_108 : _GEN_107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_110 = ~io_inputBit | _GEN_109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_111 = i == 10'h8d ? _GEN_110 : _GEN_109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_112 = io_inputBit ? 1'h0 : _GEN_111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_113 = i == 10'h8d ? _GEN_112 : _GEN_111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_114 = ~io_inputBit ? 1'h0 : _GEN_113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_115 = i == 10'h8e ? _GEN_114 : _GEN_113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_116 = io_inputBit | _GEN_115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_117 = i == 10'h8e ? _GEN_116 : _GEN_115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_118 = ~io_inputBit | _GEN_117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_119 = i == 10'h8f ? _GEN_118 : _GEN_117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_120 = io_inputBit ? 1'h0 : _GEN_119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_121 = i == 10'h8f ? _GEN_120 : _GEN_119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_122 = ~io_inputBit ? 1'h0 : _GEN_121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_123 = i == 10'h91 ? _GEN_122 : _GEN_121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_124 = io_inputBit | _GEN_123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_125 = i == 10'h91 ? _GEN_124 : _GEN_123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_126 = ~io_inputBit | _GEN_125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_127 = i == 10'h92 ? _GEN_126 : _GEN_125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_128 = io_inputBit ? 1'h0 : _GEN_127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_129 = i == 10'h92 ? _GEN_128 : _GEN_127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_130 = io_inputBit ? 1'h0 : buffer_4; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_131 = i == 10'h0 ? _GEN_130 : buffer_4; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_132 = io_inputBit ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_133 = i == 10'h1 ? _GEN_132 : _GEN_131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_134 = ~io_inputBit | _GEN_133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_135 = i == 10'h7 ? _GEN_134 : _GEN_133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_136 = io_inputBit ? 1'h0 : _GEN_135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_137 = i == 10'h8 ? _GEN_136 : _GEN_135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_138 = io_inputBit ? 1'h0 : _GEN_137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_139 = i == 10'h11 ? _GEN_138 : _GEN_137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_140 = ~io_inputBit | _GEN_139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_141 = i == 10'h21 ? _GEN_140 : _GEN_139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_142 = ~io_inputBit | _GEN_141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_143 = i == 10'h44 ? _GEN_142 : _GEN_141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_144 = ~io_inputBit ? 1'h0 : _GEN_143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_145 = i == 10'h45 ? _GEN_144 : _GEN_143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_146 = ~io_inputBit | _GEN_145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_147 = i == 10'h46 ? _GEN_146 : _GEN_145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_148 = ~io_inputBit ? 1'h0 : _GEN_147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_149 = i == 10'h47 ? _GEN_148 : _GEN_147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_150 = ~io_inputBit | _GEN_149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_151 = i == 10'h48 ? _GEN_150 : _GEN_149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_152 = ~io_inputBit ? 1'h0 : _GEN_151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_153 = i == 10'h8a ? _GEN_152 : _GEN_151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_154 = io_inputBit | _GEN_153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_155 = i == 10'h8a ? _GEN_154 : _GEN_153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_156 = ~io_inputBit | _GEN_155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_157 = i == 10'h8c ? _GEN_156 : _GEN_155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_158 = io_inputBit ? 1'h0 : _GEN_157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_159 = i == 10'h8c ? _GEN_158 : _GEN_157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_160 = ~io_inputBit ? 1'h0 : _GEN_159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_161 = i == 10'h8e ? _GEN_160 : _GEN_159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_162 = io_inputBit | _GEN_161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_163 = i == 10'h8e ? _GEN_162 : _GEN_161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_164 = ~io_inputBit | _GEN_163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_165 = i == 10'h90 ? _GEN_164 : _GEN_163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_166 = io_inputBit ? 1'h0 : _GEN_165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_167 = i == 10'h90 ? _GEN_166 : _GEN_165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_168 = ~io_inputBit ? 1'h0 : _GEN_167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_169 = i == 10'h92 ? _GEN_168 : _GEN_167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_170 = io_inputBit | _GEN_169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_171 = i == 10'h92 ? _GEN_170 : _GEN_169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_172 = io_inputBit ? 1'h0 : buffer_5; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_173 = i == 10'h0 ? _GEN_172 : buffer_5; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_174 = io_inputBit ? 1'h0 : _GEN_173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_175 = i == 10'h1 ? _GEN_174 : _GEN_173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_176 = ~io_inputBit ? 1'h0 : _GEN_175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_177 = i == 10'h7 ? _GEN_176 : _GEN_175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_178 = io_inputBit ? 1'h0 : _GEN_177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_179 = i == 10'h8 ? _GEN_178 : _GEN_177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_180 = io_inputBit ? 1'h0 : _GEN_179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_181 = i == 10'h11 ? _GEN_180 : _GEN_179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_182 = ~io_inputBit ? 1'h0 : _GEN_181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_183 = i == 10'h21 ? _GEN_182 : _GEN_181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_184 = ~io_inputBit ? 1'h0 : _GEN_183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_185 = i == 10'h89 ? _GEN_184 : _GEN_183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_186 = io_inputBit | _GEN_185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_187 = i == 10'h89 ? _GEN_186 : _GEN_185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_188 = ~io_inputBit | _GEN_187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_189 = i == 10'h8a ? _GEN_188 : _GEN_187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_190 = io_inputBit ? 1'h0 : _GEN_189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_191 = i == 10'h8a ? _GEN_190 : _GEN_189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_192 = ~io_inputBit ? 1'h0 : _GEN_191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_193 = i == 10'h8b ? _GEN_192 : _GEN_191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_194 = io_inputBit | _GEN_193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_195 = i == 10'h8b ? _GEN_194 : _GEN_193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_196 = ~io_inputBit | _GEN_195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_197 = i == 10'h8c ? _GEN_196 : _GEN_195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_198 = io_inputBit ? 1'h0 : _GEN_197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_199 = i == 10'h8c ? _GEN_198 : _GEN_197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_200 = ~io_inputBit ? 1'h0 : _GEN_199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_201 = i == 10'h8d ? _GEN_200 : _GEN_199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_202 = io_inputBit | _GEN_201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_203 = i == 10'h8d ? _GEN_202 : _GEN_201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_204 = ~io_inputBit | _GEN_203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_205 = i == 10'h8e ? _GEN_204 : _GEN_203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_206 = io_inputBit ? 1'h0 : _GEN_205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_207 = i == 10'h8e ? _GEN_206 : _GEN_205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_208 = ~io_inputBit ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_209 = i == 10'h8f ? _GEN_208 : _GEN_207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_210 = io_inputBit | _GEN_209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_211 = i == 10'h8f ? _GEN_210 : _GEN_209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_212 = ~io_inputBit | _GEN_211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_213 = i == 10'h90 ? _GEN_212 : _GEN_211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_214 = io_inputBit ? 1'h0 : _GEN_213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_215 = i == 10'h90 ? _GEN_214 : _GEN_213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_216 = ~io_inputBit ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_217 = i == 10'h91 ? _GEN_216 : _GEN_215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_218 = io_inputBit | _GEN_217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_219 = i == 10'h91 ? _GEN_218 : _GEN_217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_220 = ~io_inputBit | _GEN_219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_221 = i == 10'h92 ? _GEN_220 : _GEN_219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_222 = io_inputBit ? 1'h0 : _GEN_221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_223 = i == 10'h92 ? _GEN_222 : _GEN_221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_224 = io_inputBit ? 1'h0 : buffer_6; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_225 = i == 10'h0 ? _GEN_224 : buffer_6; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_226 = io_inputBit ? 1'h0 : _GEN_225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_227 = i == 10'h1 ? _GEN_226 : _GEN_225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_228 = ~io_inputBit ? 1'h0 : _GEN_227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_229 = i == 10'h7 ? _GEN_228 : _GEN_227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_230 = io_inputBit ? 1'h0 : _GEN_229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_231 = i == 10'h8 ? _GEN_230 : _GEN_229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_232 = io_inputBit ? 1'h0 : _GEN_231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_233 = i == 10'h11 ? _GEN_232 : _GEN_231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_234 = ~io_inputBit ? 1'h0 : _GEN_233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_235 = i == 10'h21 ? _GEN_234 : _GEN_233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_236 = ~io_inputBit ? 1'h0 : _GEN_235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_237 = i == 10'h89 ? _GEN_236 : _GEN_235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_238 = io_inputBit | _GEN_237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_239 = i == 10'h89 ? _GEN_238 : _GEN_237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_240 = ~io_inputBit ? 1'h0 : _GEN_239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_241 = i == 10'h8a ? _GEN_240 : _GEN_239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_242 = io_inputBit | _GEN_241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_243 = i == 10'h8a ? _GEN_242 : _GEN_241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_244 = ~io_inputBit ? 1'h0 : _GEN_243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_245 = i == 10'h8b ? _GEN_244 : _GEN_243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_246 = io_inputBit | _GEN_245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_247 = i == 10'h8b ? _GEN_246 : _GEN_245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_248 = ~io_inputBit ? 1'h0 : _GEN_247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_249 = i == 10'h8c ? _GEN_248 : _GEN_247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_250 = io_inputBit | _GEN_249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_251 = i == 10'h8c ? _GEN_250 : _GEN_249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_252 = ~io_inputBit ? 1'h0 : _GEN_251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_253 = i == 10'h8d ? _GEN_252 : _GEN_251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_254 = io_inputBit | _GEN_253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_255 = i == 10'h8d ? _GEN_254 : _GEN_253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_256 = ~io_inputBit ? 1'h0 : _GEN_255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_257 = i == 10'h8e ? _GEN_256 : _GEN_255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_258 = io_inputBit | _GEN_257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_259 = i == 10'h8e ? _GEN_258 : _GEN_257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_260 = ~io_inputBit ? 1'h0 : _GEN_259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_261 = i == 10'h8f ? _GEN_260 : _GEN_259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_262 = io_inputBit | _GEN_261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_263 = i == 10'h8f ? _GEN_262 : _GEN_261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_264 = ~io_inputBit ? 1'h0 : _GEN_263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_265 = i == 10'h90 ? _GEN_264 : _GEN_263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_266 = io_inputBit | _GEN_265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_267 = i == 10'h90 ? _GEN_266 : _GEN_265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_268 = ~io_inputBit ? 1'h0 : _GEN_267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_269 = i == 10'h91 ? _GEN_268 : _GEN_267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_270 = io_inputBit | _GEN_269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_271 = i == 10'h91 ? _GEN_270 : _GEN_269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_272 = ~io_inputBit ? 1'h0 : _GEN_271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_273 = i == 10'h92 ? _GEN_272 : _GEN_271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_274 = io_inputBit | _GEN_273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_275 = i == 10'h92 ? _GEN_274 : _GEN_273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_276 = io_inputBit ? 1'h0 : _GEN_13; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_277 = i == 10'h0 ? _GEN_276 : _GEN_13; // @[lut_mem_online.scala 234:34]
  wire  _GEN_278 = ~io_inputBit ? 1'h0 : _GEN_277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_279 = i == 10'h3 ? _GEN_278 : _GEN_277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_280 = io_inputBit ? 1'h0 : _GEN_279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_281 = i == 10'h4 ? _GEN_280 : _GEN_279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_282 = io_inputBit | _GEN_281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_283 = i == 10'h8 ? _GEN_282 : _GEN_281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_284 = io_inputBit ? 1'h0 : _GEN_283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_285 = i == 10'h9 ? _GEN_284 : _GEN_283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_286 = io_inputBit | _GEN_285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_287 = i == 10'h11 ? _GEN_286 : _GEN_285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_288 = io_inputBit ? 1'h0 : _GEN_287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_289 = i == 10'h13 ? _GEN_288 : _GEN_287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_290 = io_inputBit | _GEN_289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_291 = i == 10'h23 ? _GEN_290 : _GEN_289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_292 = ~io_inputBit | _GEN_291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_293 = i == 10'h27 ? _GEN_292 : _GEN_291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_294 = io_inputBit ? 1'h0 : _GEN_293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_295 = i == 10'h27 ? _GEN_294 : _GEN_293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_296 = io_inputBit | _GEN_295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_297 = i == 10'h47 ? _GEN_296 : _GEN_295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_298 = ~io_inputBit ? 1'h0 : _GEN_297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_299 = i == 10'h8f ? _GEN_298 : _GEN_297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_300 = io_inputBit | _GEN_299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_301 = i == 10'h8f ? _GEN_300 : _GEN_299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_302 = io_inputBit ? 1'h0 : _GEN_41; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_303 = i == 10'h0 ? _GEN_302 : _GEN_41; // @[lut_mem_online.scala 234:34]
  wire  _GEN_304 = io_inputBit ? 1'h0 : _GEN_303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_305 = i == 10'h4 ? _GEN_304 : _GEN_303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_306 = ~io_inputBit ? 1'h0 : _GEN_305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_307 = i == 10'h7 ? _GEN_306 : _GEN_305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_308 = io_inputBit ? 1'h0 : _GEN_307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_309 = i == 10'h9 ? _GEN_308 : _GEN_307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_310 = ~io_inputBit ? 1'h0 : _GEN_309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_311 = i == 10'h10 ? _GEN_310 : _GEN_309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_312 = io_inputBit | _GEN_311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_313 = i == 10'h11 ? _GEN_312 : _GEN_311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_314 = ~io_inputBit | _GEN_313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_315 = i == 10'h12 ? _GEN_314 : _GEN_313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_316 = io_inputBit | _GEN_315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_317 = i == 10'h22 ? _GEN_316 : _GEN_315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_318 = io_inputBit ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_319 = i == 10'h23 ? _GEN_318 : _GEN_317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_320 = ~io_inputBit | _GEN_319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_321 = i == 10'h26 ? _GEN_320 : _GEN_319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_322 = ~io_inputBit ? 1'h0 : _GEN_321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_323 = i == 10'h27 ? _GEN_322 : _GEN_321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_324 = io_inputBit | _GEN_323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_325 = i == 10'h27 ? _GEN_324 : _GEN_323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_326 = io_inputBit ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_327 = i == 10'h28 ? _GEN_326 : _GEN_325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_328 = ~io_inputBit ? 1'h0 : _GEN_327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_329 = i == 10'h45 ? _GEN_328 : _GEN_327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_330 = io_inputBit ? 1'h0 : _GEN_329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_331 = i == 10'h47 ? _GEN_330 : _GEN_329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_332 = io_inputBit ? 1'h0 : _GEN_331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_333 = i == 10'h4e ? _GEN_332 : _GEN_331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_334 = ~io_inputBit | _GEN_333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_335 = i == 10'h51 ? _GEN_334 : _GEN_333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_336 = io_inputBit ? 1'h0 : _GEN_335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_337 = i == 10'h51 ? _GEN_336 : _GEN_335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_338 = ~io_inputBit ? 1'h0 : _GEN_337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_339 = i == 10'h8c ? _GEN_338 : _GEN_337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_340 = io_inputBit | _GEN_339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_341 = i == 10'h8c ? _GEN_340 : _GEN_339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_342 = ~io_inputBit | _GEN_341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_343 = i == 10'h8f ? _GEN_342 : _GEN_341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_344 = io_inputBit ? 1'h0 : _GEN_343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_345 = i == 10'h8f ? _GEN_344 : _GEN_343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_346 = ~io_inputBit | _GEN_345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_347 = i == 10'h9d ? _GEN_346 : _GEN_345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_348 = io_inputBit ? 1'h0 : _GEN_347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_349 = i == 10'h9d ? _GEN_348 : _GEN_347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_350 = io_inputBit ? 1'h0 : _GEN_81; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_351 = i == 10'h0 ? _GEN_350 : _GEN_81; // @[lut_mem_online.scala 234:34]
  wire  _GEN_352 = io_inputBit ? 1'h0 : _GEN_351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_353 = i == 10'h4 ? _GEN_352 : _GEN_351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_354 = ~io_inputBit ? 1'h0 : _GEN_353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_355 = i == 10'h7 ? _GEN_354 : _GEN_353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_356 = io_inputBit ? 1'h0 : _GEN_355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_357 = i == 10'h9 ? _GEN_356 : _GEN_355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_358 = ~io_inputBit ? 1'h0 : _GEN_357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_359 = i == 10'h10 ? _GEN_358 : _GEN_357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_360 = io_inputBit ? 1'h0 : _GEN_359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_361 = i == 10'h11 ? _GEN_360 : _GEN_359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_362 = ~io_inputBit ? 1'h0 : _GEN_361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_363 = i == 10'h12 ? _GEN_362 : _GEN_361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_364 = io_inputBit | _GEN_363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_365 = i == 10'h23 ? _GEN_364 : _GEN_363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_366 = ~io_inputBit ? 1'h0 : _GEN_365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_367 = i == 10'h26 ? _GEN_366 : _GEN_365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_368 = ~io_inputBit | _GEN_367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_369 = i == 10'h45 ? _GEN_368 : _GEN_367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_370 = ~io_inputBit ? 1'h0 : _GEN_369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_371 = i == 10'h46 ? _GEN_370 : _GEN_369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_372 = io_inputBit | _GEN_371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_373 = i == 10'h46 ? _GEN_372 : _GEN_371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_374 = io_inputBit ? 1'h0 : _GEN_373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_375 = i == 10'h47 ? _GEN_374 : _GEN_373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_376 = io_inputBit | _GEN_375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_377 = i == 10'h4e ? _GEN_376 : _GEN_375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_378 = io_inputBit ? 1'h0 : _GEN_377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_379 = i == 10'h4f ? _GEN_378 : _GEN_377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_380 = ~io_inputBit | _GEN_379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_381 = i == 10'h50 ? _GEN_380 : _GEN_379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_382 = ~io_inputBit ? 1'h0 : _GEN_381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_383 = i == 10'h51 ? _GEN_382 : _GEN_381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_384 = io_inputBit | _GEN_383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_385 = i == 10'h51 ? _GEN_384 : _GEN_383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_386 = io_inputBit ? 1'h0 : _GEN_385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_387 = i == 10'h52 ? _GEN_386 : _GEN_385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_388 = ~io_inputBit | _GEN_387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_389 = i == 10'h8c ? _GEN_388 : _GEN_387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_390 = io_inputBit ? 1'h0 : _GEN_389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_391 = i == 10'h8c ? _GEN_390 : _GEN_389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_392 = ~io_inputBit | _GEN_391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_393 = i == 10'h8f ? _GEN_392 : _GEN_391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_394 = io_inputBit ? 1'h0 : _GEN_393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_395 = i == 10'h8f ? _GEN_394 : _GEN_393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_396 = ~io_inputBit ? 1'h0 : _GEN_395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_397 = i == 10'h9d ? _GEN_396 : _GEN_395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_398 = io_inputBit | _GEN_397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_399 = i == 10'h9d ? _GEN_398 : _GEN_397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_400 = ~io_inputBit | _GEN_399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_401 = i == 10'h9f ? _GEN_400 : _GEN_399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_402 = io_inputBit ? 1'h0 : _GEN_401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_403 = i == 10'h9f ? _GEN_402 : _GEN_401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_404 = ~io_inputBit | _GEN_403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_405 = i == 10'ha2 ? _GEN_404 : _GEN_403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_406 = io_inputBit ? 1'h0 : _GEN_405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_407 = i == 10'ha2 ? _GEN_406 : _GEN_405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_408 = ~io_inputBit | _GEN_407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_409 = i == 10'ha5 ? _GEN_408 : _GEN_407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_410 = io_inputBit ? 1'h0 : _GEN_409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_411 = i == 10'ha5 ? _GEN_410 : _GEN_409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_412 = io_inputBit ? 1'h0 : _GEN_129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_413 = i == 10'h0 ? _GEN_412 : _GEN_129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_414 = io_inputBit ? 1'h0 : _GEN_413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_415 = i == 10'h4 ? _GEN_414 : _GEN_413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_416 = ~io_inputBit ? 1'h0 : _GEN_415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_417 = i == 10'h7 ? _GEN_416 : _GEN_415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_418 = io_inputBit ? 1'h0 : _GEN_417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_419 = i == 10'h9 ? _GEN_418 : _GEN_417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_420 = io_inputBit ? 1'h0 : _GEN_419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_421 = i == 10'h11 ? _GEN_420 : _GEN_419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_422 = ~io_inputBit ? 1'h0 : _GEN_421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_423 = i == 10'h12 ? _GEN_422 : _GEN_421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_424 = ~io_inputBit ? 1'h0 : _GEN_423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_425 = i == 10'h21 ? _GEN_424 : _GEN_423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_426 = ~io_inputBit ? 1'h0 : _GEN_425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_427 = i == 10'h26 ? _GEN_426 : _GEN_425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_428 = ~io_inputBit ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_429 = i == 10'h44 ? _GEN_428 : _GEN_427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_430 = io_inputBit | _GEN_429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_431 = i == 10'h44 ? _GEN_430 : _GEN_429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_432 = ~io_inputBit | _GEN_431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_433 = i == 10'h46 ? _GEN_432 : _GEN_431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_434 = io_inputBit ? 1'h0 : _GEN_433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_435 = i == 10'h46 ? _GEN_434 : _GEN_433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_436 = ~io_inputBit ? 1'h0 : _GEN_435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_437 = i == 10'h48 ? _GEN_436 : _GEN_435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_438 = io_inputBit | _GEN_437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_439 = i == 10'h48 ? _GEN_438 : _GEN_437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_440 = io_inputBit ? 1'h0 : _GEN_439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_441 = i == 10'h4f ? _GEN_440 : _GEN_439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_442 = io_inputBit | _GEN_441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_443 = i == 10'h51 ? _GEN_442 : _GEN_441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_444 = ~io_inputBit ? 1'h0 : _GEN_443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_445 = i == 10'h8b ? _GEN_444 : _GEN_443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_446 = io_inputBit | _GEN_445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_447 = i == 10'h8b ? _GEN_446 : _GEN_445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_448 = ~io_inputBit | _GEN_447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_449 = i == 10'h8c ? _GEN_448 : _GEN_447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_450 = io_inputBit ? 1'h0 : _GEN_449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_451 = i == 10'h8c ? _GEN_450 : _GEN_449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_452 = ~io_inputBit | _GEN_451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_453 = i == 10'h8f ? _GEN_452 : _GEN_451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_454 = io_inputBit ? 1'h0 : _GEN_453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_455 = i == 10'h8f ? _GEN_454 : _GEN_453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_456 = ~io_inputBit ? 1'h0 : _GEN_455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_457 = i == 10'h90 ? _GEN_456 : _GEN_455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_458 = io_inputBit | _GEN_457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_459 = i == 10'h90 ? _GEN_458 : _GEN_457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_460 = ~io_inputBit ? 1'h0 : _GEN_459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_461 = i == 10'h9d ? _GEN_460 : _GEN_459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_462 = io_inputBit | _GEN_461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_463 = i == 10'h9d ? _GEN_462 : _GEN_461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_464 = ~io_inputBit | _GEN_463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_465 = i == 10'h9e ? _GEN_464 : _GEN_463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_466 = io_inputBit ? 1'h0 : _GEN_465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_467 = i == 10'h9e ? _GEN_466 : _GEN_465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_468 = ~io_inputBit ? 1'h0 : _GEN_467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_469 = i == 10'h9f ? _GEN_468 : _GEN_467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_470 = io_inputBit | _GEN_469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_471 = i == 10'h9f ? _GEN_470 : _GEN_469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_472 = ~io_inputBit | _GEN_471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_473 = i == 10'ha1 ? _GEN_472 : _GEN_471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_474 = io_inputBit ? 1'h0 : _GEN_473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_475 = i == 10'ha1 ? _GEN_474 : _GEN_473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_476 = ~io_inputBit ? 1'h0 : _GEN_475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_477 = i == 10'ha2 ? _GEN_476 : _GEN_475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_478 = io_inputBit | _GEN_477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_479 = i == 10'ha2 ? _GEN_478 : _GEN_477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_480 = ~io_inputBit | _GEN_479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_481 = i == 10'ha3 ? _GEN_480 : _GEN_479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_482 = io_inputBit ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_483 = i == 10'ha3 ? _GEN_482 : _GEN_481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_484 = ~io_inputBit ? 1'h0 : _GEN_483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_485 = i == 10'ha5 ? _GEN_484 : _GEN_483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_486 = io_inputBit | _GEN_485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_487 = i == 10'ha5 ? _GEN_486 : _GEN_485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_488 = ~io_inputBit | _GEN_487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_489 = i == 10'ha6 ? _GEN_488 : _GEN_487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_490 = io_inputBit ? 1'h0 : _GEN_489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_491 = i == 10'ha6 ? _GEN_490 : _GEN_489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_492 = io_inputBit ? 1'h0 : _GEN_171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_493 = i == 10'h0 ? _GEN_492 : _GEN_171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_494 = io_inputBit ? 1'h0 : _GEN_493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_495 = i == 10'h4 ? _GEN_494 : _GEN_493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_496 = ~io_inputBit ? 1'h0 : _GEN_495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_497 = i == 10'h7 ? _GEN_496 : _GEN_495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_498 = io_inputBit ? 1'h0 : _GEN_497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_499 = i == 10'h9 ? _GEN_498 : _GEN_497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_500 = io_inputBit | _GEN_499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_501 = i == 10'h11 ? _GEN_500 : _GEN_499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_502 = ~io_inputBit | _GEN_501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_503 = i == 10'h12 ? _GEN_502 : _GEN_501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_504 = ~io_inputBit ? 1'h0 : _GEN_503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_505 = i == 10'h21 ? _GEN_504 : _GEN_503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_506 = ~io_inputBit | _GEN_505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_507 = i == 10'h26 ? _GEN_506 : _GEN_505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_508 = ~io_inputBit | _GEN_507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_509 = i == 10'h4e ? _GEN_508 : _GEN_507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_510 = ~io_inputBit ? 1'h0 : _GEN_509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_511 = i == 10'h4f ? _GEN_510 : _GEN_509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_512 = ~io_inputBit | _GEN_511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_513 = i == 10'h50 ? _GEN_512 : _GEN_511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_514 = ~io_inputBit ? 1'h0 : _GEN_513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_515 = i == 10'h51 ? _GEN_514 : _GEN_513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_516 = ~io_inputBit | _GEN_515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_517 = i == 10'h52 ? _GEN_516 : _GEN_515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_518 = ~io_inputBit ? 1'h0 : _GEN_517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_519 = i == 10'h89 ? _GEN_518 : _GEN_517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_520 = io_inputBit | _GEN_519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_521 = i == 10'h89 ? _GEN_520 : _GEN_519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_522 = ~io_inputBit ? 1'h0 : _GEN_521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_523 = i == 10'h8a ? _GEN_522 : _GEN_521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_524 = io_inputBit | _GEN_523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_525 = i == 10'h8a ? _GEN_524 : _GEN_523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_526 = ~io_inputBit | _GEN_525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_527 = i == 10'h8b ? _GEN_526 : _GEN_525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_528 = io_inputBit ? 1'h0 : _GEN_527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_529 = i == 10'h8b ? _GEN_528 : _GEN_527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_530 = ~io_inputBit | _GEN_529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_531 = i == 10'h8c ? _GEN_530 : _GEN_529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_532 = io_inputBit ? 1'h0 : _GEN_531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_533 = i == 10'h8c ? _GEN_532 : _GEN_531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_534 = ~io_inputBit ? 1'h0 : _GEN_533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_535 = i == 10'h8d ? _GEN_534 : _GEN_533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_536 = io_inputBit | _GEN_535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_537 = i == 10'h8d ? _GEN_536 : _GEN_535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_538 = ~io_inputBit ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_539 = i == 10'h8e ? _GEN_538 : _GEN_537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_540 = io_inputBit | _GEN_539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_541 = i == 10'h8e ? _GEN_540 : _GEN_539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_542 = ~io_inputBit | _GEN_541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_543 = i == 10'h8f ? _GEN_542 : _GEN_541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_544 = io_inputBit ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_545 = i == 10'h8f ? _GEN_544 : _GEN_543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_546 = ~io_inputBit | _GEN_545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_547 = i == 10'h90 ? _GEN_546 : _GEN_545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_548 = io_inputBit ? 1'h0 : _GEN_547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_549 = i == 10'h90 ? _GEN_548 : _GEN_547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_550 = ~io_inputBit ? 1'h0 : _GEN_549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_551 = i == 10'h91 ? _GEN_550 : _GEN_549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_552 = io_inputBit | _GEN_551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_553 = i == 10'h91 ? _GEN_552 : _GEN_551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_554 = ~io_inputBit ? 1'h0 : _GEN_553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_555 = i == 10'h92 ? _GEN_554 : _GEN_553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_556 = io_inputBit | _GEN_555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_557 = i == 10'h92 ? _GEN_556 : _GEN_555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_558 = ~io_inputBit ? 1'h0 : _GEN_557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_559 = i == 10'h9e ? _GEN_558 : _GEN_557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_560 = io_inputBit | _GEN_559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_561 = i == 10'h9e ? _GEN_560 : _GEN_559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_562 = ~io_inputBit | _GEN_561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_563 = i == 10'ha0 ? _GEN_562 : _GEN_561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_564 = io_inputBit ? 1'h0 : _GEN_563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_565 = i == 10'ha0 ? _GEN_564 : _GEN_563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_566 = ~io_inputBit ? 1'h0 : _GEN_565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_567 = i == 10'ha2 ? _GEN_566 : _GEN_565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_568 = io_inputBit | _GEN_567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_569 = i == 10'ha2 ? _GEN_568 : _GEN_567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_570 = ~io_inputBit | _GEN_569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_571 = i == 10'ha4 ? _GEN_570 : _GEN_569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_572 = io_inputBit ? 1'h0 : _GEN_571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_573 = i == 10'ha4 ? _GEN_572 : _GEN_571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_574 = ~io_inputBit ? 1'h0 : _GEN_573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_575 = i == 10'ha6 ? _GEN_574 : _GEN_573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_576 = io_inputBit | _GEN_575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_577 = i == 10'ha6 ? _GEN_576 : _GEN_575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_578 = io_inputBit ? 1'h0 : _GEN_223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_579 = i == 10'h0 ? _GEN_578 : _GEN_223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_580 = io_inputBit ? 1'h0 : _GEN_579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_581 = i == 10'h4 ? _GEN_580 : _GEN_579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_582 = ~io_inputBit ? 1'h0 : _GEN_581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_583 = i == 10'h7 ? _GEN_582 : _GEN_581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_584 = io_inputBit ? 1'h0 : _GEN_583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_585 = i == 10'h9 ? _GEN_584 : _GEN_583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_586 = io_inputBit ? 1'h0 : _GEN_585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_587 = i == 10'h11 ? _GEN_586 : _GEN_585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_588 = ~io_inputBit ? 1'h0 : _GEN_587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_589 = i == 10'h12 ? _GEN_588 : _GEN_587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_590 = ~io_inputBit ? 1'h0 : _GEN_589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_591 = i == 10'h21 ? _GEN_590 : _GEN_589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_592 = ~io_inputBit ? 1'h0 : _GEN_591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_593 = i == 10'h26 ? _GEN_592 : _GEN_591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_594 = ~io_inputBit ? 1'h0 : _GEN_593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_595 = i == 10'h44 ? _GEN_594 : _GEN_593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_596 = io_inputBit | _GEN_595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_597 = i == 10'h44 ? _GEN_596 : _GEN_595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_598 = ~io_inputBit ? 1'h0 : _GEN_597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_599 = i == 10'h45 ? _GEN_598 : _GEN_597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_600 = io_inputBit | _GEN_599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_601 = i == 10'h45 ? _GEN_600 : _GEN_599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_602 = ~io_inputBit ? 1'h0 : _GEN_601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_603 = i == 10'h46 ? _GEN_602 : _GEN_601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_604 = io_inputBit | _GEN_603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_605 = i == 10'h46 ? _GEN_604 : _GEN_603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_606 = ~io_inputBit ? 1'h0 : _GEN_605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_607 = i == 10'h47 ? _GEN_606 : _GEN_605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_608 = io_inputBit | _GEN_607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_609 = i == 10'h47 ? _GEN_608 : _GEN_607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_610 = ~io_inputBit ? 1'h0 : _GEN_609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_611 = i == 10'h48 ? _GEN_610 : _GEN_609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_612 = io_inputBit | _GEN_611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_613 = i == 10'h48 ? _GEN_612 : _GEN_611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_614 = ~io_inputBit ? 1'h0 : _GEN_613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_615 = i == 10'h9d ? _GEN_614 : _GEN_613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_616 = io_inputBit | _GEN_615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_617 = i == 10'h9d ? _GEN_616 : _GEN_615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_618 = ~io_inputBit | _GEN_617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_619 = i == 10'h9e ? _GEN_618 : _GEN_617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_620 = io_inputBit ? 1'h0 : _GEN_619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_621 = i == 10'h9e ? _GEN_620 : _GEN_619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_622 = ~io_inputBit ? 1'h0 : _GEN_621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_623 = i == 10'h9f ? _GEN_622 : _GEN_621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_624 = io_inputBit | _GEN_623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_625 = i == 10'h9f ? _GEN_624 : _GEN_623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_626 = ~io_inputBit | _GEN_625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_627 = i == 10'ha0 ? _GEN_626 : _GEN_625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_628 = io_inputBit ? 1'h0 : _GEN_627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_629 = i == 10'ha0 ? _GEN_628 : _GEN_627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_630 = ~io_inputBit ? 1'h0 : _GEN_629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_631 = i == 10'ha1 ? _GEN_630 : _GEN_629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_632 = io_inputBit | _GEN_631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_633 = i == 10'ha1 ? _GEN_632 : _GEN_631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_634 = ~io_inputBit | _GEN_633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_635 = i == 10'ha2 ? _GEN_634 : _GEN_633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_636 = io_inputBit ? 1'h0 : _GEN_635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_637 = i == 10'ha2 ? _GEN_636 : _GEN_635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_638 = ~io_inputBit ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_639 = i == 10'ha3 ? _GEN_638 : _GEN_637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_640 = io_inputBit | _GEN_639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_641 = i == 10'ha3 ? _GEN_640 : _GEN_639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_642 = ~io_inputBit | _GEN_641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_643 = i == 10'ha4 ? _GEN_642 : _GEN_641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_644 = io_inputBit ? 1'h0 : _GEN_643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_645 = i == 10'ha4 ? _GEN_644 : _GEN_643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_646 = ~io_inputBit ? 1'h0 : _GEN_645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_647 = i == 10'ha5 ? _GEN_646 : _GEN_645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_648 = io_inputBit | _GEN_647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_649 = i == 10'ha5 ? _GEN_648 : _GEN_647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_650 = ~io_inputBit | _GEN_649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_651 = i == 10'ha6 ? _GEN_650 : _GEN_649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_652 = io_inputBit ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_653 = i == 10'ha6 ? _GEN_652 : _GEN_651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_654 = io_inputBit ? 1'h0 : _GEN_275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_655 = i == 10'h0 ? _GEN_654 : _GEN_275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_656 = io_inputBit ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_657 = i == 10'h4 ? _GEN_656 : _GEN_655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_658 = ~io_inputBit ? 1'h0 : _GEN_657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_659 = i == 10'h7 ? _GEN_658 : _GEN_657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_660 = io_inputBit ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_661 = i == 10'h9 ? _GEN_660 : _GEN_659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_662 = io_inputBit ? 1'h0 : _GEN_661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_663 = i == 10'h11 ? _GEN_662 : _GEN_661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_664 = ~io_inputBit ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_665 = i == 10'h12 ? _GEN_664 : _GEN_663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_666 = ~io_inputBit ? 1'h0 : _GEN_665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_667 = i == 10'h21 ? _GEN_666 : _GEN_665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_668 = ~io_inputBit ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_669 = i == 10'h26 ? _GEN_668 : _GEN_667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_670 = ~io_inputBit ? 1'h0 : _GEN_669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_671 = i == 10'h89 ? _GEN_670 : _GEN_669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_672 = io_inputBit | _GEN_671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_673 = i == 10'h89 ? _GEN_672 : _GEN_671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_674 = ~io_inputBit ? 1'h0 : _GEN_673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_675 = i == 10'h8a ? _GEN_674 : _GEN_673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_676 = io_inputBit | _GEN_675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_677 = i == 10'h8a ? _GEN_676 : _GEN_675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_678 = ~io_inputBit ? 1'h0 : _GEN_677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_679 = i == 10'h8b ? _GEN_678 : _GEN_677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_680 = io_inputBit | _GEN_679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_681 = i == 10'h8b ? _GEN_680 : _GEN_679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_682 = ~io_inputBit ? 1'h0 : _GEN_681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_683 = i == 10'h8c ? _GEN_682 : _GEN_681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_684 = io_inputBit | _GEN_683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_685 = i == 10'h8c ? _GEN_684 : _GEN_683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_686 = ~io_inputBit ? 1'h0 : _GEN_685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_687 = i == 10'h8d ? _GEN_686 : _GEN_685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_688 = io_inputBit | _GEN_687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_689 = i == 10'h8d ? _GEN_688 : _GEN_687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_690 = ~io_inputBit ? 1'h0 : _GEN_689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_691 = i == 10'h8e ? _GEN_690 : _GEN_689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_692 = io_inputBit | _GEN_691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_693 = i == 10'h8e ? _GEN_692 : _GEN_691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_694 = ~io_inputBit ? 1'h0 : _GEN_693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_695 = i == 10'h8f ? _GEN_694 : _GEN_693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_696 = io_inputBit | _GEN_695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_697 = i == 10'h8f ? _GEN_696 : _GEN_695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_698 = ~io_inputBit ? 1'h0 : _GEN_697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_699 = i == 10'h90 ? _GEN_698 : _GEN_697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_700 = io_inputBit | _GEN_699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_701 = i == 10'h90 ? _GEN_700 : _GEN_699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_702 = ~io_inputBit ? 1'h0 : _GEN_701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_703 = i == 10'h91 ? _GEN_702 : _GEN_701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_704 = io_inputBit | _GEN_703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_705 = i == 10'h91 ? _GEN_704 : _GEN_703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_706 = ~io_inputBit ? 1'h0 : _GEN_705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_707 = i == 10'h92 ? _GEN_706 : _GEN_705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_708 = io_inputBit | _GEN_707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_709 = i == 10'h92 ? _GEN_708 : _GEN_707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_710 = ~io_inputBit ? 1'h0 : _GEN_709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_711 = i == 10'h9d ? _GEN_710 : _GEN_709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_712 = io_inputBit | _GEN_711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_713 = i == 10'h9d ? _GEN_712 : _GEN_711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_714 = ~io_inputBit ? 1'h0 : _GEN_713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_715 = i == 10'h9e ? _GEN_714 : _GEN_713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_716 = io_inputBit | _GEN_715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_717 = i == 10'h9e ? _GEN_716 : _GEN_715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_718 = ~io_inputBit ? 1'h0 : _GEN_717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_719 = i == 10'h9f ? _GEN_718 : _GEN_717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_720 = io_inputBit | _GEN_719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_721 = i == 10'h9f ? _GEN_720 : _GEN_719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_722 = ~io_inputBit ? 1'h0 : _GEN_721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_723 = i == 10'ha0 ? _GEN_722 : _GEN_721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_724 = io_inputBit | _GEN_723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_725 = i == 10'ha0 ? _GEN_724 : _GEN_723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_726 = ~io_inputBit ? 1'h0 : _GEN_725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_727 = i == 10'ha1 ? _GEN_726 : _GEN_725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_728 = io_inputBit | _GEN_727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_729 = i == 10'ha1 ? _GEN_728 : _GEN_727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_730 = ~io_inputBit ? 1'h0 : _GEN_729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_731 = i == 10'ha2 ? _GEN_730 : _GEN_729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_732 = io_inputBit | _GEN_731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_733 = i == 10'ha2 ? _GEN_732 : _GEN_731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_734 = ~io_inputBit ? 1'h0 : _GEN_733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_735 = i == 10'ha3 ? _GEN_734 : _GEN_733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_736 = io_inputBit | _GEN_735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_737 = i == 10'ha3 ? _GEN_736 : _GEN_735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_738 = ~io_inputBit ? 1'h0 : _GEN_737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_739 = i == 10'ha4 ? _GEN_738 : _GEN_737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_740 = io_inputBit | _GEN_739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_741 = i == 10'ha4 ? _GEN_740 : _GEN_739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_742 = ~io_inputBit ? 1'h0 : _GEN_741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_743 = i == 10'ha5 ? _GEN_742 : _GEN_741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_744 = io_inputBit | _GEN_743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_745 = i == 10'ha5 ? _GEN_744 : _GEN_743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_746 = ~io_inputBit ? 1'h0 : _GEN_745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_747 = i == 10'ha6 ? _GEN_746 : _GEN_745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_748 = io_inputBit | _GEN_747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_749 = i == 10'ha6 ? _GEN_748 : _GEN_747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_750 = io_inputBit ? 1'h0 : _GEN_301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_751 = i == 10'h0 ? _GEN_750 : _GEN_301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_752 = ~io_inputBit ? 1'h0 : _GEN_751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_753 = i == 10'h1 ? _GEN_752 : _GEN_751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_754 = io_inputBit | _GEN_753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_755 = i == 10'h9 ? _GEN_754 : _GEN_753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_756 = io_inputBit ? 1'h0 : _GEN_755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_757 = i == 10'ha ? _GEN_756 : _GEN_755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_758 = ~io_inputBit ? 1'h0 : _GEN_757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_759 = i == 10'h13 ? _GEN_758 : _GEN_757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_760 = ~io_inputBit | _GEN_759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_761 = i == 10'h15 ? _GEN_760 : _GEN_759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_762 = io_inputBit | _GEN_761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_763 = i == 10'h28 ? _GEN_762 : _GEN_761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_764 = ~io_inputBit | _GEN_763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_765 = i == 10'h2c ? _GEN_764 : _GEN_763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_766 = io_inputBit ? 1'h0 : _GEN_765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_767 = i == 10'h2c ? _GEN_766 : _GEN_765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_768 = io_inputBit | _GEN_767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_769 = i == 10'h51 ? _GEN_768 : _GEN_767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_770 = ~io_inputBit ? 1'h0 : _GEN_769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_771 = i == 10'ha3 ? _GEN_770 : _GEN_769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_772 = io_inputBit | _GEN_771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_773 = i == 10'ha3 ? _GEN_772 : _GEN_771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_774 = io_inputBit ? 1'h0 : _GEN_349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_775 = i == 10'h0 ? _GEN_774 : _GEN_349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_776 = ~io_inputBit ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_777 = i == 10'h1 ? _GEN_776 : _GEN_775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_778 = io_inputBit | _GEN_777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_779 = i == 10'h9 ? _GEN_778 : _GEN_777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_780 = io_inputBit ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_781 = i == 10'h16 ? _GEN_780 : _GEN_779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_782 = io_inputBit | _GEN_781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_783 = i == 10'h27 ? _GEN_782 : _GEN_781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_784 = io_inputBit ? 1'h0 : _GEN_783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_785 = i == 10'h28 ? _GEN_784 : _GEN_783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_786 = ~io_inputBit | _GEN_785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_787 = i == 10'h2b ? _GEN_786 : _GEN_785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_788 = ~io_inputBit ? 1'h0 : _GEN_787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_789 = i == 10'h2c ? _GEN_788 : _GEN_787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_790 = io_inputBit | _GEN_789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_791 = i == 10'h2c ? _GEN_790 : _GEN_789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_792 = io_inputBit ? 1'h0 : _GEN_791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_793 = i == 10'h2d ? _GEN_792 : _GEN_791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_794 = ~io_inputBit ? 1'h0 : _GEN_793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_795 = i == 10'h4f ? _GEN_794 : _GEN_793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_796 = io_inputBit ? 1'h0 : _GEN_795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_797 = i == 10'h51 ? _GEN_796 : _GEN_795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_798 = io_inputBit ? 1'h0 : _GEN_797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_799 = i == 10'h58 ? _GEN_798 : _GEN_797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_800 = ~io_inputBit | _GEN_799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_801 = i == 10'h5b ? _GEN_800 : _GEN_799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_802 = io_inputBit ? 1'h0 : _GEN_801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_803 = i == 10'h5b ? _GEN_802 : _GEN_801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_804 = ~io_inputBit ? 1'h0 : _GEN_803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_805 = i == 10'ha0 ? _GEN_804 : _GEN_803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_806 = io_inputBit | _GEN_805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_807 = i == 10'ha0 ? _GEN_806 : _GEN_805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_808 = ~io_inputBit | _GEN_807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_809 = i == 10'ha3 ? _GEN_808 : _GEN_807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_810 = io_inputBit ? 1'h0 : _GEN_809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_811 = i == 10'ha3 ? _GEN_810 : _GEN_809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_812 = ~io_inputBit | _GEN_811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_813 = i == 10'hb1 ? _GEN_812 : _GEN_811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_814 = io_inputBit ? 1'h0 : _GEN_813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_815 = i == 10'hb1 ? _GEN_814 : _GEN_813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_816 = io_inputBit ? 1'h0 : _GEN_411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_817 = i == 10'h0 ? _GEN_816 : _GEN_411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_818 = ~io_inputBit ? 1'h0 : _GEN_817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_819 = i == 10'h1 ? _GEN_818 : _GEN_817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_820 = io_inputBit ? 1'h0 : _GEN_819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_821 = i == 10'h9 ? _GEN_820 : _GEN_819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_822 = io_inputBit ? 1'h0 : _GEN_821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_823 = i == 10'h16 ? _GEN_822 : _GEN_821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_824 = io_inputBit | _GEN_823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_825 = i == 10'h28 ? _GEN_824 : _GEN_823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_826 = ~io_inputBit ? 1'h0 : _GEN_825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_827 = i == 10'h2b ? _GEN_826 : _GEN_825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_828 = ~io_inputBit | _GEN_827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_829 = i == 10'h4f ? _GEN_828 : _GEN_827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_830 = ~io_inputBit ? 1'h0 : _GEN_829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_831 = i == 10'h50 ? _GEN_830 : _GEN_829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_832 = io_inputBit | _GEN_831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_833 = i == 10'h50 ? _GEN_832 : _GEN_831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_834 = io_inputBit ? 1'h0 : _GEN_833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_835 = i == 10'h51 ? _GEN_834 : _GEN_833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_836 = io_inputBit | _GEN_835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_837 = i == 10'h58 ? _GEN_836 : _GEN_835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_838 = io_inputBit ? 1'h0 : _GEN_837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_839 = i == 10'h59 ? _GEN_838 : _GEN_837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_840 = ~io_inputBit | _GEN_839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_841 = i == 10'h5a ? _GEN_840 : _GEN_839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_842 = ~io_inputBit ? 1'h0 : _GEN_841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_843 = i == 10'h5b ? _GEN_842 : _GEN_841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_844 = io_inputBit | _GEN_843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_845 = i == 10'h5b ? _GEN_844 : _GEN_843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_846 = io_inputBit ? 1'h0 : _GEN_845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_847 = i == 10'h5c ? _GEN_846 : _GEN_845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_848 = ~io_inputBit | _GEN_847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_849 = i == 10'ha0 ? _GEN_848 : _GEN_847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_850 = io_inputBit ? 1'h0 : _GEN_849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_851 = i == 10'ha0 ? _GEN_850 : _GEN_849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_852 = ~io_inputBit | _GEN_851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_853 = i == 10'ha3 ? _GEN_852 : _GEN_851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_854 = io_inputBit ? 1'h0 : _GEN_853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_855 = i == 10'ha3 ? _GEN_854 : _GEN_853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_856 = ~io_inputBit ? 1'h0 : _GEN_855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_857 = i == 10'hb1 ? _GEN_856 : _GEN_855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_858 = io_inputBit | _GEN_857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_859 = i == 10'hb1 ? _GEN_858 : _GEN_857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_860 = ~io_inputBit | _GEN_859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_861 = i == 10'hb3 ? _GEN_860 : _GEN_859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_862 = io_inputBit ? 1'h0 : _GEN_861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_863 = i == 10'hb3 ? _GEN_862 : _GEN_861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_864 = ~io_inputBit | _GEN_863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_865 = i == 10'hb6 ? _GEN_864 : _GEN_863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_866 = io_inputBit ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_867 = i == 10'hb6 ? _GEN_866 : _GEN_865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_868 = ~io_inputBit | _GEN_867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_869 = i == 10'hb9 ? _GEN_868 : _GEN_867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_870 = io_inputBit ? 1'h0 : _GEN_869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_871 = i == 10'hb9 ? _GEN_870 : _GEN_869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_872 = io_inputBit ? 1'h0 : _GEN_491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_873 = i == 10'h0 ? _GEN_872 : _GEN_491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_874 = ~io_inputBit ? 1'h0 : _GEN_873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_875 = i == 10'h3 ? _GEN_874 : _GEN_873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_876 = ~io_inputBit ? 1'h0 : _GEN_875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_877 = i == 10'h8 ? _GEN_876 : _GEN_875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_878 = io_inputBit ? 1'h0 : _GEN_877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_879 = i == 10'h9 ? _GEN_878 : _GEN_877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_880 = ~io_inputBit ? 1'h0 : _GEN_879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_881 = i == 10'h12 ? _GEN_880 : _GEN_879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_882 = io_inputBit ? 1'h0 : _GEN_881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_883 = i == 10'h16 ? _GEN_882 : _GEN_881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_884 = ~io_inputBit ? 1'h0 : _GEN_883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_885 = i == 10'h26 ? _GEN_884 : _GEN_883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_886 = ~io_inputBit ? 1'h0 : _GEN_885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_887 = i == 10'h2b ? _GEN_886 : _GEN_885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_888 = ~io_inputBit ? 1'h0 : _GEN_887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_889 = i == 10'h4e ? _GEN_888 : _GEN_887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_890 = io_inputBit | _GEN_889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_891 = i == 10'h4e ? _GEN_890 : _GEN_889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_892 = ~io_inputBit | _GEN_891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_893 = i == 10'h50 ? _GEN_892 : _GEN_891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_894 = io_inputBit ? 1'h0 : _GEN_893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_895 = i == 10'h50 ? _GEN_894 : _GEN_893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_896 = ~io_inputBit ? 1'h0 : _GEN_895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_897 = i == 10'h52 ? _GEN_896 : _GEN_895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_898 = io_inputBit | _GEN_897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_899 = i == 10'h52 ? _GEN_898 : _GEN_897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_900 = io_inputBit ? 1'h0 : _GEN_899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_901 = i == 10'h59 ? _GEN_900 : _GEN_899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_902 = io_inputBit | _GEN_901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_903 = i == 10'h5b ? _GEN_902 : _GEN_901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_904 = ~io_inputBit ? 1'h0 : _GEN_903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_905 = i == 10'h9f ? _GEN_904 : _GEN_903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_906 = io_inputBit | _GEN_905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_907 = i == 10'h9f ? _GEN_906 : _GEN_905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_908 = ~io_inputBit | _GEN_907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_909 = i == 10'ha0 ? _GEN_908 : _GEN_907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_910 = io_inputBit ? 1'h0 : _GEN_909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_911 = i == 10'ha0 ? _GEN_910 : _GEN_909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_912 = ~io_inputBit | _GEN_911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_913 = i == 10'ha3 ? _GEN_912 : _GEN_911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_914 = io_inputBit ? 1'h0 : _GEN_913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_915 = i == 10'ha3 ? _GEN_914 : _GEN_913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_916 = ~io_inputBit ? 1'h0 : _GEN_915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_917 = i == 10'ha4 ? _GEN_916 : _GEN_915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_918 = io_inputBit | _GEN_917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_919 = i == 10'ha4 ? _GEN_918 : _GEN_917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_920 = ~io_inputBit ? 1'h0 : _GEN_919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_921 = i == 10'hb1 ? _GEN_920 : _GEN_919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_922 = io_inputBit | _GEN_921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_923 = i == 10'hb1 ? _GEN_922 : _GEN_921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_924 = ~io_inputBit | _GEN_923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_925 = i == 10'hb2 ? _GEN_924 : _GEN_923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_926 = io_inputBit ? 1'h0 : _GEN_925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_927 = i == 10'hb2 ? _GEN_926 : _GEN_925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_928 = ~io_inputBit ? 1'h0 : _GEN_927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_929 = i == 10'hb3 ? _GEN_928 : _GEN_927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_930 = io_inputBit | _GEN_929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_931 = i == 10'hb3 ? _GEN_930 : _GEN_929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_932 = ~io_inputBit | _GEN_931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_933 = i == 10'hb5 ? _GEN_932 : _GEN_931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_934 = io_inputBit ? 1'h0 : _GEN_933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_935 = i == 10'hb5 ? _GEN_934 : _GEN_933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_936 = ~io_inputBit ? 1'h0 : _GEN_935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_937 = i == 10'hb6 ? _GEN_936 : _GEN_935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_938 = io_inputBit | _GEN_937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_939 = i == 10'hb6 ? _GEN_938 : _GEN_937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_940 = ~io_inputBit | _GEN_939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_941 = i == 10'hb7 ? _GEN_940 : _GEN_939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_942 = io_inputBit ? 1'h0 : _GEN_941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_943 = i == 10'hb7 ? _GEN_942 : _GEN_941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_944 = ~io_inputBit ? 1'h0 : _GEN_943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_945 = i == 10'hb9 ? _GEN_944 : _GEN_943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_946 = io_inputBit | _GEN_945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_947 = i == 10'hb9 ? _GEN_946 : _GEN_945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_948 = ~io_inputBit | _GEN_947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_949 = i == 10'hba ? _GEN_948 : _GEN_947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_950 = io_inputBit ? 1'h0 : _GEN_949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_951 = i == 10'hba ? _GEN_950 : _GEN_949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_952 = io_inputBit ? 1'h0 : _GEN_577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_953 = i == 10'h0 ? _GEN_952 : _GEN_577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_954 = ~io_inputBit ? 1'h0 : _GEN_953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_955 = i == 10'h3 ? _GEN_954 : _GEN_953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_956 = ~io_inputBit ? 1'h0 : _GEN_955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_957 = i == 10'h8 ? _GEN_956 : _GEN_955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_958 = io_inputBit | _GEN_957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_959 = i == 10'h9 ? _GEN_958 : _GEN_957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_960 = ~io_inputBit ? 1'h0 : _GEN_959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_961 = i == 10'h12 ? _GEN_960 : _GEN_959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_962 = io_inputBit ? 1'h0 : _GEN_961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_963 = i == 10'h16 ? _GEN_962 : _GEN_961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_964 = ~io_inputBit ? 1'h0 : _GEN_963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_965 = i == 10'h26 ? _GEN_964 : _GEN_963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_966 = ~io_inputBit | _GEN_965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_967 = i == 10'h2b ? _GEN_966 : _GEN_965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_968 = ~io_inputBit | _GEN_967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_969 = i == 10'h58 ? _GEN_968 : _GEN_967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_970 = ~io_inputBit ? 1'h0 : _GEN_969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_971 = i == 10'h59 ? _GEN_970 : _GEN_969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_972 = ~io_inputBit | _GEN_971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_973 = i == 10'h5a ? _GEN_972 : _GEN_971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_974 = ~io_inputBit ? 1'h0 : _GEN_973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_975 = i == 10'h5b ? _GEN_974 : _GEN_973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_976 = ~io_inputBit | _GEN_975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_977 = i == 10'h5c ? _GEN_976 : _GEN_975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_978 = ~io_inputBit ? 1'h0 : _GEN_977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_979 = i == 10'h9d ? _GEN_978 : _GEN_977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_980 = io_inputBit | _GEN_979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_981 = i == 10'h9d ? _GEN_980 : _GEN_979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_982 = ~io_inputBit ? 1'h0 : _GEN_981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_983 = i == 10'h9e ? _GEN_982 : _GEN_981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_984 = io_inputBit | _GEN_983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_985 = i == 10'h9e ? _GEN_984 : _GEN_983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_986 = ~io_inputBit | _GEN_985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_987 = i == 10'h9f ? _GEN_986 : _GEN_985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_988 = io_inputBit ? 1'h0 : _GEN_987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_989 = i == 10'h9f ? _GEN_988 : _GEN_987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_990 = ~io_inputBit | _GEN_989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_991 = i == 10'ha0 ? _GEN_990 : _GEN_989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_992 = io_inputBit ? 1'h0 : _GEN_991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_993 = i == 10'ha0 ? _GEN_992 : _GEN_991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_994 = ~io_inputBit ? 1'h0 : _GEN_993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_995 = i == 10'ha1 ? _GEN_994 : _GEN_993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_996 = io_inputBit | _GEN_995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_997 = i == 10'ha1 ? _GEN_996 : _GEN_995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_998 = ~io_inputBit ? 1'h0 : _GEN_997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_999 = i == 10'ha2 ? _GEN_998 : _GEN_997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1000 = io_inputBit | _GEN_999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1001 = i == 10'ha2 ? _GEN_1000 : _GEN_999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1002 = ~io_inputBit | _GEN_1001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1003 = i == 10'ha3 ? _GEN_1002 : _GEN_1001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1004 = io_inputBit ? 1'h0 : _GEN_1003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1005 = i == 10'ha3 ? _GEN_1004 : _GEN_1003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1006 = ~io_inputBit | _GEN_1005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1007 = i == 10'ha4 ? _GEN_1006 : _GEN_1005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1008 = io_inputBit ? 1'h0 : _GEN_1007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1009 = i == 10'ha4 ? _GEN_1008 : _GEN_1007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1010 = ~io_inputBit ? 1'h0 : _GEN_1009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1011 = i == 10'ha5 ? _GEN_1010 : _GEN_1009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1012 = io_inputBit | _GEN_1011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1013 = i == 10'ha5 ? _GEN_1012 : _GEN_1011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1014 = ~io_inputBit ? 1'h0 : _GEN_1013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1015 = i == 10'ha6 ? _GEN_1014 : _GEN_1013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1016 = io_inputBit | _GEN_1015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1017 = i == 10'ha6 ? _GEN_1016 : _GEN_1015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1018 = ~io_inputBit ? 1'h0 : _GEN_1017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1019 = i == 10'hb2 ? _GEN_1018 : _GEN_1017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1020 = io_inputBit | _GEN_1019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1021 = i == 10'hb2 ? _GEN_1020 : _GEN_1019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1022 = ~io_inputBit | _GEN_1021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1023 = i == 10'hb4 ? _GEN_1022 : _GEN_1021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1024 = io_inputBit ? 1'h0 : _GEN_1023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1025 = i == 10'hb4 ? _GEN_1024 : _GEN_1023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1026 = ~io_inputBit ? 1'h0 : _GEN_1025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1027 = i == 10'hb6 ? _GEN_1026 : _GEN_1025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1028 = io_inputBit | _GEN_1027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1029 = i == 10'hb6 ? _GEN_1028 : _GEN_1027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1030 = ~io_inputBit | _GEN_1029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1031 = i == 10'hb8 ? _GEN_1030 : _GEN_1029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1032 = io_inputBit ? 1'h0 : _GEN_1031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1033 = i == 10'hb8 ? _GEN_1032 : _GEN_1031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1034 = ~io_inputBit ? 1'h0 : _GEN_1033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1035 = i == 10'hba ? _GEN_1034 : _GEN_1033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1036 = io_inputBit | _GEN_1035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1037 = i == 10'hba ? _GEN_1036 : _GEN_1035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1038 = io_inputBit ? 1'h0 : _GEN_653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1039 = i == 10'h0 ? _GEN_1038 : _GEN_653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1040 = ~io_inputBit ? 1'h0 : _GEN_1039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1041 = i == 10'h3 ? _GEN_1040 : _GEN_1039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1042 = ~io_inputBit ? 1'h0 : _GEN_1041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1043 = i == 10'h8 ? _GEN_1042 : _GEN_1041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1044 = io_inputBit ? 1'h0 : _GEN_1043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1045 = i == 10'h9 ? _GEN_1044 : _GEN_1043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1046 = ~io_inputBit ? 1'h0 : _GEN_1045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1047 = i == 10'h12 ? _GEN_1046 : _GEN_1045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1048 = io_inputBit ? 1'h0 : _GEN_1047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1049 = i == 10'h16 ? _GEN_1048 : _GEN_1047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1050 = ~io_inputBit ? 1'h0 : _GEN_1049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1051 = i == 10'h26 ? _GEN_1050 : _GEN_1049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1052 = ~io_inputBit ? 1'h0 : _GEN_1051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1053 = i == 10'h2b ? _GEN_1052 : _GEN_1051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1054 = ~io_inputBit ? 1'h0 : _GEN_1053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1055 = i == 10'h4e ? _GEN_1054 : _GEN_1053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1056 = io_inputBit | _GEN_1055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1057 = i == 10'h4e ? _GEN_1056 : _GEN_1055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1058 = ~io_inputBit ? 1'h0 : _GEN_1057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1059 = i == 10'h4f ? _GEN_1058 : _GEN_1057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1060 = io_inputBit | _GEN_1059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1061 = i == 10'h4f ? _GEN_1060 : _GEN_1059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1062 = ~io_inputBit ? 1'h0 : _GEN_1061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1063 = i == 10'h50 ? _GEN_1062 : _GEN_1061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1064 = io_inputBit | _GEN_1063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1065 = i == 10'h50 ? _GEN_1064 : _GEN_1063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1066 = ~io_inputBit ? 1'h0 : _GEN_1065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1067 = i == 10'h51 ? _GEN_1066 : _GEN_1065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1068 = io_inputBit | _GEN_1067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1069 = i == 10'h51 ? _GEN_1068 : _GEN_1067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1070 = ~io_inputBit ? 1'h0 : _GEN_1069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1071 = i == 10'h52 ? _GEN_1070 : _GEN_1069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1072 = io_inputBit | _GEN_1071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1073 = i == 10'h52 ? _GEN_1072 : _GEN_1071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1074 = ~io_inputBit ? 1'h0 : _GEN_1073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1075 = i == 10'hb1 ? _GEN_1074 : _GEN_1073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1076 = io_inputBit | _GEN_1075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1077 = i == 10'hb1 ? _GEN_1076 : _GEN_1075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1078 = ~io_inputBit | _GEN_1077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1079 = i == 10'hb2 ? _GEN_1078 : _GEN_1077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1080 = io_inputBit ? 1'h0 : _GEN_1079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1081 = i == 10'hb2 ? _GEN_1080 : _GEN_1079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1082 = ~io_inputBit ? 1'h0 : _GEN_1081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1083 = i == 10'hb3 ? _GEN_1082 : _GEN_1081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1084 = io_inputBit | _GEN_1083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1085 = i == 10'hb3 ? _GEN_1084 : _GEN_1083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1086 = ~io_inputBit | _GEN_1085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1087 = i == 10'hb4 ? _GEN_1086 : _GEN_1085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1088 = io_inputBit ? 1'h0 : _GEN_1087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1089 = i == 10'hb4 ? _GEN_1088 : _GEN_1087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1090 = ~io_inputBit ? 1'h0 : _GEN_1089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1091 = i == 10'hb5 ? _GEN_1090 : _GEN_1089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1092 = io_inputBit | _GEN_1091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1093 = i == 10'hb5 ? _GEN_1092 : _GEN_1091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1094 = ~io_inputBit | _GEN_1093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1095 = i == 10'hb6 ? _GEN_1094 : _GEN_1093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1096 = io_inputBit ? 1'h0 : _GEN_1095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1097 = i == 10'hb6 ? _GEN_1096 : _GEN_1095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1098 = ~io_inputBit ? 1'h0 : _GEN_1097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1099 = i == 10'hb7 ? _GEN_1098 : _GEN_1097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1100 = io_inputBit | _GEN_1099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1101 = i == 10'hb7 ? _GEN_1100 : _GEN_1099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1102 = ~io_inputBit | _GEN_1101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1103 = i == 10'hb8 ? _GEN_1102 : _GEN_1101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1104 = io_inputBit ? 1'h0 : _GEN_1103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1105 = i == 10'hb8 ? _GEN_1104 : _GEN_1103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1106 = ~io_inputBit ? 1'h0 : _GEN_1105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1107 = i == 10'hb9 ? _GEN_1106 : _GEN_1105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1108 = io_inputBit | _GEN_1107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1109 = i == 10'hb9 ? _GEN_1108 : _GEN_1107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1110 = ~io_inputBit | _GEN_1109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1111 = i == 10'hba ? _GEN_1110 : _GEN_1109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1112 = io_inputBit ? 1'h0 : _GEN_1111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1113 = i == 10'hba ? _GEN_1112 : _GEN_1111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1114 = io_inputBit ? 1'h0 : _GEN_749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1115 = i == 10'h0 ? _GEN_1114 : _GEN_749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1116 = ~io_inputBit ? 1'h0 : _GEN_1115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1117 = i == 10'h3 ? _GEN_1116 : _GEN_1115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1118 = ~io_inputBit ? 1'h0 : _GEN_1117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1119 = i == 10'h8 ? _GEN_1118 : _GEN_1117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1120 = io_inputBit ? 1'h0 : _GEN_1119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1121 = i == 10'h9 ? _GEN_1120 : _GEN_1119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1122 = ~io_inputBit ? 1'h0 : _GEN_1121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1123 = i == 10'h12 ? _GEN_1122 : _GEN_1121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1124 = io_inputBit ? 1'h0 : _GEN_1123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1125 = i == 10'h16 ? _GEN_1124 : _GEN_1123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1126 = ~io_inputBit ? 1'h0 : _GEN_1125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1127 = i == 10'h26 ? _GEN_1126 : _GEN_1125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1128 = ~io_inputBit ? 1'h0 : _GEN_1127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1129 = i == 10'h2b ? _GEN_1128 : _GEN_1127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1130 = ~io_inputBit ? 1'h0 : _GEN_1129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1131 = i == 10'h9d ? _GEN_1130 : _GEN_1129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1132 = io_inputBit | _GEN_1131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1133 = i == 10'h9d ? _GEN_1132 : _GEN_1131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1134 = ~io_inputBit ? 1'h0 : _GEN_1133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1135 = i == 10'h9e ? _GEN_1134 : _GEN_1133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1136 = io_inputBit | _GEN_1135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1137 = i == 10'h9e ? _GEN_1136 : _GEN_1135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1138 = ~io_inputBit ? 1'h0 : _GEN_1137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1139 = i == 10'h9f ? _GEN_1138 : _GEN_1137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1140 = io_inputBit | _GEN_1139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1141 = i == 10'h9f ? _GEN_1140 : _GEN_1139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1142 = ~io_inputBit ? 1'h0 : _GEN_1141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1143 = i == 10'ha0 ? _GEN_1142 : _GEN_1141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1144 = io_inputBit | _GEN_1143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1145 = i == 10'ha0 ? _GEN_1144 : _GEN_1143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1146 = ~io_inputBit ? 1'h0 : _GEN_1145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1147 = i == 10'ha1 ? _GEN_1146 : _GEN_1145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1148 = io_inputBit | _GEN_1147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1149 = i == 10'ha1 ? _GEN_1148 : _GEN_1147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1150 = ~io_inputBit ? 1'h0 : _GEN_1149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1151 = i == 10'ha2 ? _GEN_1150 : _GEN_1149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1152 = io_inputBit | _GEN_1151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1153 = i == 10'ha2 ? _GEN_1152 : _GEN_1151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1154 = ~io_inputBit ? 1'h0 : _GEN_1153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1155 = i == 10'ha3 ? _GEN_1154 : _GEN_1153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1156 = io_inputBit | _GEN_1155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1157 = i == 10'ha3 ? _GEN_1156 : _GEN_1155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1158 = ~io_inputBit ? 1'h0 : _GEN_1157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1159 = i == 10'ha4 ? _GEN_1158 : _GEN_1157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1160 = io_inputBit | _GEN_1159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1161 = i == 10'ha4 ? _GEN_1160 : _GEN_1159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1162 = ~io_inputBit ? 1'h0 : _GEN_1161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1163 = i == 10'ha5 ? _GEN_1162 : _GEN_1161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1164 = io_inputBit | _GEN_1163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1165 = i == 10'ha5 ? _GEN_1164 : _GEN_1163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1166 = ~io_inputBit ? 1'h0 : _GEN_1165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1167 = i == 10'ha6 ? _GEN_1166 : _GEN_1165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1168 = io_inputBit | _GEN_1167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1169 = i == 10'ha6 ? _GEN_1168 : _GEN_1167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1170 = ~io_inputBit ? 1'h0 : _GEN_1169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1171 = i == 10'hb1 ? _GEN_1170 : _GEN_1169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1172 = io_inputBit | _GEN_1171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1173 = i == 10'hb1 ? _GEN_1172 : _GEN_1171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1174 = ~io_inputBit ? 1'h0 : _GEN_1173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1175 = i == 10'hb2 ? _GEN_1174 : _GEN_1173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1176 = io_inputBit | _GEN_1175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1177 = i == 10'hb2 ? _GEN_1176 : _GEN_1175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1178 = ~io_inputBit ? 1'h0 : _GEN_1177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1179 = i == 10'hb3 ? _GEN_1178 : _GEN_1177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1180 = io_inputBit | _GEN_1179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1181 = i == 10'hb3 ? _GEN_1180 : _GEN_1179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1182 = ~io_inputBit ? 1'h0 : _GEN_1181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1183 = i == 10'hb4 ? _GEN_1182 : _GEN_1181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1184 = io_inputBit | _GEN_1183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1185 = i == 10'hb4 ? _GEN_1184 : _GEN_1183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1186 = ~io_inputBit ? 1'h0 : _GEN_1185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1187 = i == 10'hb5 ? _GEN_1186 : _GEN_1185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1188 = io_inputBit | _GEN_1187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1189 = i == 10'hb5 ? _GEN_1188 : _GEN_1187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1190 = ~io_inputBit ? 1'h0 : _GEN_1189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1191 = i == 10'hb6 ? _GEN_1190 : _GEN_1189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1192 = io_inputBit | _GEN_1191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1193 = i == 10'hb6 ? _GEN_1192 : _GEN_1191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1194 = ~io_inputBit ? 1'h0 : _GEN_1193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1195 = i == 10'hb7 ? _GEN_1194 : _GEN_1193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1196 = io_inputBit | _GEN_1195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1197 = i == 10'hb7 ? _GEN_1196 : _GEN_1195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1198 = ~io_inputBit ? 1'h0 : _GEN_1197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1199 = i == 10'hb8 ? _GEN_1198 : _GEN_1197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1200 = io_inputBit | _GEN_1199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1201 = i == 10'hb8 ? _GEN_1200 : _GEN_1199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1202 = ~io_inputBit ? 1'h0 : _GEN_1201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1203 = i == 10'hb9 ? _GEN_1202 : _GEN_1201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1204 = io_inputBit | _GEN_1203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1205 = i == 10'hb9 ? _GEN_1204 : _GEN_1203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1206 = ~io_inputBit ? 1'h0 : _GEN_1205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1207 = i == 10'hba ? _GEN_1206 : _GEN_1205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1208 = io_inputBit | _GEN_1207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1209 = i == 10'hba ? _GEN_1208 : _GEN_1207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1210 = ~io_inputBit ? 1'h0 : _GEN_773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1211 = i == 10'h1 ? _GEN_1210 : _GEN_773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1212 = io_inputBit ? 1'h0 : _GEN_1211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1213 = i == 10'h2 ? _GEN_1212 : _GEN_1211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1214 = ~io_inputBit ? 1'h0 : _GEN_1213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1215 = i == 10'h4 ? _GEN_1214 : _GEN_1213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1216 = io_inputBit ? 1'h0 : _GEN_1215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1217 = i == 10'h5 ? _GEN_1216 : _GEN_1215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1218 = ~io_inputBit ? 1'h0 : _GEN_1217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1219 = i == 10'ha ? _GEN_1218 : _GEN_1217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1220 = ~io_inputBit | _GEN_1219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1221 = i == 10'hb ? _GEN_1220 : _GEN_1219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1222 = io_inputBit | _GEN_1221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1223 = i == 10'h16 ? _GEN_1222 : _GEN_1221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1224 = io_inputBit ? 1'h0 : _GEN_1223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1225 = i == 10'h18 ? _GEN_1224 : _GEN_1223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1226 = io_inputBit | _GEN_1225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1227 = i == 10'h2d ? _GEN_1226 : _GEN_1225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1228 = ~io_inputBit | _GEN_1227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1229 = i == 10'h31 ? _GEN_1228 : _GEN_1227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1230 = io_inputBit ? 1'h0 : _GEN_1229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1231 = i == 10'h31 ? _GEN_1230 : _GEN_1229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1232 = io_inputBit | _GEN_1231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1233 = i == 10'h5b ? _GEN_1232 : _GEN_1231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1234 = ~io_inputBit ? 1'h0 : _GEN_1233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1235 = i == 10'hb7 ? _GEN_1234 : _GEN_1233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1236 = io_inputBit | _GEN_1235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1237 = i == 10'hb7 ? _GEN_1236 : _GEN_1235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1238 = ~io_inputBit ? 1'h0 : _GEN_815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1239 = i == 10'h1 ? _GEN_1238 : _GEN_815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1240 = io_inputBit ? 1'h0 : _GEN_1239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1241 = i == 10'h2 ? _GEN_1240 : _GEN_1239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1242 = ~io_inputBit ? 1'h0 : _GEN_1241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1243 = i == 10'h4 ? _GEN_1242 : _GEN_1241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1244 = io_inputBit ? 1'h0 : _GEN_1243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1245 = i == 10'h5 ? _GEN_1244 : _GEN_1243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1246 = ~io_inputBit ? 1'h0 : _GEN_1245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1247 = i == 10'h15 ? _GEN_1246 : _GEN_1245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1248 = io_inputBit | _GEN_1247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1249 = i == 10'h16 ? _GEN_1248 : _GEN_1247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1250 = ~io_inputBit | _GEN_1249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1251 = i == 10'h17 ? _GEN_1250 : _GEN_1249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1252 = io_inputBit | _GEN_1251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1253 = i == 10'h2c ? _GEN_1252 : _GEN_1251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1254 = io_inputBit ? 1'h0 : _GEN_1253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1255 = i == 10'h2d ? _GEN_1254 : _GEN_1253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1256 = ~io_inputBit | _GEN_1255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1257 = i == 10'h30 ? _GEN_1256 : _GEN_1255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1258 = ~io_inputBit ? 1'h0 : _GEN_1257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1259 = i == 10'h31 ? _GEN_1258 : _GEN_1257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1260 = io_inputBit | _GEN_1259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1261 = i == 10'h31 ? _GEN_1260 : _GEN_1259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1262 = io_inputBit ? 1'h0 : _GEN_1261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1263 = i == 10'h32 ? _GEN_1262 : _GEN_1261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1264 = ~io_inputBit ? 1'h0 : _GEN_1263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1265 = i == 10'h59 ? _GEN_1264 : _GEN_1263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1266 = io_inputBit ? 1'h0 : _GEN_1265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1267 = i == 10'h5b ? _GEN_1266 : _GEN_1265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1268 = io_inputBit ? 1'h0 : _GEN_1267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1269 = i == 10'h62 ? _GEN_1268 : _GEN_1267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1270 = ~io_inputBit | _GEN_1269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1271 = i == 10'h65 ? _GEN_1270 : _GEN_1269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1272 = io_inputBit ? 1'h0 : _GEN_1271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1273 = i == 10'h65 ? _GEN_1272 : _GEN_1271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1274 = ~io_inputBit ? 1'h0 : _GEN_1273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1275 = i == 10'hb4 ? _GEN_1274 : _GEN_1273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1276 = io_inputBit | _GEN_1275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1277 = i == 10'hb4 ? _GEN_1276 : _GEN_1275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1278 = ~io_inputBit | _GEN_1277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1279 = i == 10'hb7 ? _GEN_1278 : _GEN_1277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1280 = io_inputBit ? 1'h0 : _GEN_1279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1281 = i == 10'hb7 ? _GEN_1280 : _GEN_1279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1282 = ~io_inputBit | _GEN_1281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1283 = i == 10'hc5 ? _GEN_1282 : _GEN_1281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1284 = io_inputBit ? 1'h0 : _GEN_1283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1285 = i == 10'hc5 ? _GEN_1284 : _GEN_1283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1286 = ~io_inputBit ? 1'h0 : _GEN_871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1287 = i == 10'h1 ? _GEN_1286 : _GEN_871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1288 = io_inputBit ? 1'h0 : _GEN_1287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1289 = i == 10'h2 ? _GEN_1288 : _GEN_1287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1290 = ~io_inputBit ? 1'h0 : _GEN_1289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1291 = i == 10'h4 ? _GEN_1290 : _GEN_1289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1292 = io_inputBit ? 1'h0 : _GEN_1291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1293 = i == 10'h5 ? _GEN_1292 : _GEN_1291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1294 = ~io_inputBit ? 1'h0 : _GEN_1293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1295 = i == 10'h15 ? _GEN_1294 : _GEN_1293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1296 = io_inputBit ? 1'h0 : _GEN_1295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1297 = i == 10'h16 ? _GEN_1296 : _GEN_1295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1298 = ~io_inputBit ? 1'h0 : _GEN_1297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1299 = i == 10'h17 ? _GEN_1298 : _GEN_1297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1300 = io_inputBit | _GEN_1299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1301 = i == 10'h2d ? _GEN_1300 : _GEN_1299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1302 = ~io_inputBit ? 1'h0 : _GEN_1301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1303 = i == 10'h30 ? _GEN_1302 : _GEN_1301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1304 = ~io_inputBit | _GEN_1303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1305 = i == 10'h59 ? _GEN_1304 : _GEN_1303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1306 = ~io_inputBit ? 1'h0 : _GEN_1305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1307 = i == 10'h5a ? _GEN_1306 : _GEN_1305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1308 = io_inputBit | _GEN_1307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1309 = i == 10'h5a ? _GEN_1308 : _GEN_1307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1310 = io_inputBit ? 1'h0 : _GEN_1309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1311 = i == 10'h5b ? _GEN_1310 : _GEN_1309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1312 = io_inputBit | _GEN_1311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1313 = i == 10'h62 ? _GEN_1312 : _GEN_1311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1314 = io_inputBit ? 1'h0 : _GEN_1313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1315 = i == 10'h63 ? _GEN_1314 : _GEN_1313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1316 = ~io_inputBit | _GEN_1315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1317 = i == 10'h64 ? _GEN_1316 : _GEN_1315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1318 = ~io_inputBit ? 1'h0 : _GEN_1317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1319 = i == 10'h65 ? _GEN_1318 : _GEN_1317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1320 = io_inputBit | _GEN_1319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1321 = i == 10'h65 ? _GEN_1320 : _GEN_1319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1322 = io_inputBit ? 1'h0 : _GEN_1321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1323 = i == 10'h66 ? _GEN_1322 : _GEN_1321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1324 = ~io_inputBit | _GEN_1323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1325 = i == 10'hb4 ? _GEN_1324 : _GEN_1323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1326 = io_inputBit ? 1'h0 : _GEN_1325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1327 = i == 10'hb4 ? _GEN_1326 : _GEN_1325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1328 = ~io_inputBit | _GEN_1327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1329 = i == 10'hb7 ? _GEN_1328 : _GEN_1327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1330 = io_inputBit ? 1'h0 : _GEN_1329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1331 = i == 10'hb7 ? _GEN_1330 : _GEN_1329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1332 = ~io_inputBit ? 1'h0 : _GEN_1331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1333 = i == 10'hc5 ? _GEN_1332 : _GEN_1331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1334 = io_inputBit | _GEN_1333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1335 = i == 10'hc5 ? _GEN_1334 : _GEN_1333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1336 = ~io_inputBit | _GEN_1335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1337 = i == 10'hc7 ? _GEN_1336 : _GEN_1335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1338 = io_inputBit ? 1'h0 : _GEN_1337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1339 = i == 10'hc7 ? _GEN_1338 : _GEN_1337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1340 = ~io_inputBit | _GEN_1339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1341 = i == 10'hca ? _GEN_1340 : _GEN_1339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1342 = io_inputBit ? 1'h0 : _GEN_1341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1343 = i == 10'hca ? _GEN_1342 : _GEN_1341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1344 = ~io_inputBit | _GEN_1343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1345 = i == 10'hcd ? _GEN_1344 : _GEN_1343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1346 = io_inputBit ? 1'h0 : _GEN_1345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1347 = i == 10'hcd ? _GEN_1346 : _GEN_1345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1348 = ~io_inputBit ? 1'h0 : _GEN_951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1349 = i == 10'h1 ? _GEN_1348 : _GEN_951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1350 = io_inputBit ? 1'h0 : _GEN_1349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1351 = i == 10'h2 ? _GEN_1350 : _GEN_1349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1352 = ~io_inputBit ? 1'h0 : _GEN_1351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1353 = i == 10'h4 ? _GEN_1352 : _GEN_1351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1354 = io_inputBit ? 1'h0 : _GEN_1353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1355 = i == 10'h5 ? _GEN_1354 : _GEN_1353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1356 = io_inputBit ? 1'h0 : _GEN_1355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1357 = i == 10'h16 ? _GEN_1356 : _GEN_1355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1358 = ~io_inputBit ? 1'h0 : _GEN_1357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1359 = i == 10'h17 ? _GEN_1358 : _GEN_1357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1360 = ~io_inputBit ? 1'h0 : _GEN_1359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1361 = i == 10'h2b ? _GEN_1360 : _GEN_1359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1362 = ~io_inputBit ? 1'h0 : _GEN_1361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1363 = i == 10'h30 ? _GEN_1362 : _GEN_1361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1364 = ~io_inputBit ? 1'h0 : _GEN_1363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1365 = i == 10'h58 ? _GEN_1364 : _GEN_1363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1366 = io_inputBit | _GEN_1365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1367 = i == 10'h58 ? _GEN_1366 : _GEN_1365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1368 = ~io_inputBit | _GEN_1367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1369 = i == 10'h5a ? _GEN_1368 : _GEN_1367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1370 = io_inputBit ? 1'h0 : _GEN_1369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1371 = i == 10'h5a ? _GEN_1370 : _GEN_1369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1372 = ~io_inputBit ? 1'h0 : _GEN_1371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1373 = i == 10'h5c ? _GEN_1372 : _GEN_1371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1374 = io_inputBit | _GEN_1373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1375 = i == 10'h5c ? _GEN_1374 : _GEN_1373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1376 = io_inputBit ? 1'h0 : _GEN_1375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1377 = i == 10'h63 ? _GEN_1376 : _GEN_1375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1378 = io_inputBit | _GEN_1377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1379 = i == 10'h65 ? _GEN_1378 : _GEN_1377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1380 = ~io_inputBit ? 1'h0 : _GEN_1379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1381 = i == 10'hb3 ? _GEN_1380 : _GEN_1379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1382 = io_inputBit | _GEN_1381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1383 = i == 10'hb3 ? _GEN_1382 : _GEN_1381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1384 = ~io_inputBit | _GEN_1383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1385 = i == 10'hb4 ? _GEN_1384 : _GEN_1383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1386 = io_inputBit ? 1'h0 : _GEN_1385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1387 = i == 10'hb4 ? _GEN_1386 : _GEN_1385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1388 = ~io_inputBit | _GEN_1387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1389 = i == 10'hb7 ? _GEN_1388 : _GEN_1387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1390 = io_inputBit ? 1'h0 : _GEN_1389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1391 = i == 10'hb7 ? _GEN_1390 : _GEN_1389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1392 = ~io_inputBit ? 1'h0 : _GEN_1391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1393 = i == 10'hb8 ? _GEN_1392 : _GEN_1391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1394 = io_inputBit | _GEN_1393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1395 = i == 10'hb8 ? _GEN_1394 : _GEN_1393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1396 = ~io_inputBit ? 1'h0 : _GEN_1395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1397 = i == 10'hc5 ? _GEN_1396 : _GEN_1395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1398 = io_inputBit | _GEN_1397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1399 = i == 10'hc5 ? _GEN_1398 : _GEN_1397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1400 = ~io_inputBit | _GEN_1399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1401 = i == 10'hc6 ? _GEN_1400 : _GEN_1399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1402 = io_inputBit ? 1'h0 : _GEN_1401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1403 = i == 10'hc6 ? _GEN_1402 : _GEN_1401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1404 = ~io_inputBit ? 1'h0 : _GEN_1403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1405 = i == 10'hc7 ? _GEN_1404 : _GEN_1403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1406 = io_inputBit | _GEN_1405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1407 = i == 10'hc7 ? _GEN_1406 : _GEN_1405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1408 = ~io_inputBit | _GEN_1407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1409 = i == 10'hc9 ? _GEN_1408 : _GEN_1407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1410 = io_inputBit ? 1'h0 : _GEN_1409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1411 = i == 10'hc9 ? _GEN_1410 : _GEN_1409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1412 = ~io_inputBit ? 1'h0 : _GEN_1411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1413 = i == 10'hca ? _GEN_1412 : _GEN_1411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1414 = io_inputBit | _GEN_1413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1415 = i == 10'hca ? _GEN_1414 : _GEN_1413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1416 = ~io_inputBit | _GEN_1415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1417 = i == 10'hcb ? _GEN_1416 : _GEN_1415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1418 = io_inputBit ? 1'h0 : _GEN_1417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1419 = i == 10'hcb ? _GEN_1418 : _GEN_1417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1420 = ~io_inputBit ? 1'h0 : _GEN_1419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1421 = i == 10'hcd ? _GEN_1420 : _GEN_1419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1422 = io_inputBit | _GEN_1421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1423 = i == 10'hcd ? _GEN_1422 : _GEN_1421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1424 = ~io_inputBit | _GEN_1423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1425 = i == 10'hce ? _GEN_1424 : _GEN_1423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1426 = io_inputBit ? 1'h0 : _GEN_1425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1427 = i == 10'hce ? _GEN_1426 : _GEN_1425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1428 = ~io_inputBit ? 1'h0 : _GEN_1037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1429 = i == 10'h1 ? _GEN_1428 : _GEN_1037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1430 = io_inputBit ? 1'h0 : _GEN_1429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1431 = i == 10'h2 ? _GEN_1430 : _GEN_1429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1432 = ~io_inputBit ? 1'h0 : _GEN_1431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1433 = i == 10'h4 ? _GEN_1432 : _GEN_1431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1434 = io_inputBit ? 1'h0 : _GEN_1433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1435 = i == 10'h5 ? _GEN_1434 : _GEN_1433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1436 = io_inputBit | _GEN_1435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1437 = i == 10'h16 ? _GEN_1436 : _GEN_1435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1438 = ~io_inputBit | _GEN_1437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1439 = i == 10'h17 ? _GEN_1438 : _GEN_1437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1440 = ~io_inputBit ? 1'h0 : _GEN_1439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1441 = i == 10'h2b ? _GEN_1440 : _GEN_1439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1442 = ~io_inputBit | _GEN_1441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1443 = i == 10'h30 ? _GEN_1442 : _GEN_1441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1444 = ~io_inputBit | _GEN_1443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1445 = i == 10'h62 ? _GEN_1444 : _GEN_1443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1446 = ~io_inputBit ? 1'h0 : _GEN_1445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1447 = i == 10'h63 ? _GEN_1446 : _GEN_1445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1448 = ~io_inputBit | _GEN_1447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1449 = i == 10'h64 ? _GEN_1448 : _GEN_1447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1450 = ~io_inputBit ? 1'h0 : _GEN_1449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1451 = i == 10'h65 ? _GEN_1450 : _GEN_1449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1452 = ~io_inputBit | _GEN_1451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1453 = i == 10'h66 ? _GEN_1452 : _GEN_1451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1454 = ~io_inputBit ? 1'h0 : _GEN_1453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1455 = i == 10'hb1 ? _GEN_1454 : _GEN_1453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1456 = io_inputBit | _GEN_1455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1457 = i == 10'hb1 ? _GEN_1456 : _GEN_1455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1458 = ~io_inputBit ? 1'h0 : _GEN_1457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1459 = i == 10'hb2 ? _GEN_1458 : _GEN_1457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1460 = io_inputBit | _GEN_1459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1461 = i == 10'hb2 ? _GEN_1460 : _GEN_1459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1462 = ~io_inputBit | _GEN_1461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1463 = i == 10'hb3 ? _GEN_1462 : _GEN_1461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1464 = io_inputBit ? 1'h0 : _GEN_1463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1465 = i == 10'hb3 ? _GEN_1464 : _GEN_1463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1466 = ~io_inputBit | _GEN_1465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1467 = i == 10'hb4 ? _GEN_1466 : _GEN_1465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1468 = io_inputBit ? 1'h0 : _GEN_1467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1469 = i == 10'hb4 ? _GEN_1468 : _GEN_1467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1470 = ~io_inputBit ? 1'h0 : _GEN_1469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1471 = i == 10'hb5 ? _GEN_1470 : _GEN_1469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1472 = io_inputBit | _GEN_1471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1473 = i == 10'hb5 ? _GEN_1472 : _GEN_1471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1474 = ~io_inputBit ? 1'h0 : _GEN_1473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1475 = i == 10'hb6 ? _GEN_1474 : _GEN_1473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1476 = io_inputBit | _GEN_1475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1477 = i == 10'hb6 ? _GEN_1476 : _GEN_1475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1478 = ~io_inputBit | _GEN_1477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1479 = i == 10'hb7 ? _GEN_1478 : _GEN_1477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1480 = io_inputBit ? 1'h0 : _GEN_1479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1481 = i == 10'hb7 ? _GEN_1480 : _GEN_1479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1482 = ~io_inputBit | _GEN_1481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1483 = i == 10'hb8 ? _GEN_1482 : _GEN_1481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1484 = io_inputBit ? 1'h0 : _GEN_1483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1485 = i == 10'hb8 ? _GEN_1484 : _GEN_1483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1486 = ~io_inputBit ? 1'h0 : _GEN_1485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1487 = i == 10'hb9 ? _GEN_1486 : _GEN_1485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1488 = io_inputBit | _GEN_1487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1489 = i == 10'hb9 ? _GEN_1488 : _GEN_1487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1490 = ~io_inputBit ? 1'h0 : _GEN_1489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1491 = i == 10'hba ? _GEN_1490 : _GEN_1489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1492 = io_inputBit | _GEN_1491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1493 = i == 10'hba ? _GEN_1492 : _GEN_1491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1494 = ~io_inputBit ? 1'h0 : _GEN_1493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1495 = i == 10'hc6 ? _GEN_1494 : _GEN_1493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1496 = io_inputBit | _GEN_1495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1497 = i == 10'hc6 ? _GEN_1496 : _GEN_1495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1498 = ~io_inputBit | _GEN_1497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1499 = i == 10'hc8 ? _GEN_1498 : _GEN_1497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1500 = io_inputBit ? 1'h0 : _GEN_1499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1501 = i == 10'hc8 ? _GEN_1500 : _GEN_1499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1502 = ~io_inputBit ? 1'h0 : _GEN_1501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1503 = i == 10'hca ? _GEN_1502 : _GEN_1501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1504 = io_inputBit | _GEN_1503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1505 = i == 10'hca ? _GEN_1504 : _GEN_1503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1506 = ~io_inputBit | _GEN_1505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1507 = i == 10'hcc ? _GEN_1506 : _GEN_1505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1508 = io_inputBit ? 1'h0 : _GEN_1507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1509 = i == 10'hcc ? _GEN_1508 : _GEN_1507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1510 = ~io_inputBit ? 1'h0 : _GEN_1509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1511 = i == 10'hce ? _GEN_1510 : _GEN_1509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1512 = io_inputBit | _GEN_1511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1513 = i == 10'hce ? _GEN_1512 : _GEN_1511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1514 = ~io_inputBit ? 1'h0 : _GEN_1113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1515 = i == 10'h1 ? _GEN_1514 : _GEN_1113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1516 = io_inputBit ? 1'h0 : _GEN_1515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1517 = i == 10'h2 ? _GEN_1516 : _GEN_1515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1518 = ~io_inputBit ? 1'h0 : _GEN_1517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1519 = i == 10'h4 ? _GEN_1518 : _GEN_1517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1520 = io_inputBit ? 1'h0 : _GEN_1519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1521 = i == 10'h5 ? _GEN_1520 : _GEN_1519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1522 = io_inputBit ? 1'h0 : _GEN_1521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1523 = i == 10'h16 ? _GEN_1522 : _GEN_1521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1524 = ~io_inputBit ? 1'h0 : _GEN_1523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1525 = i == 10'h17 ? _GEN_1524 : _GEN_1523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1526 = ~io_inputBit ? 1'h0 : _GEN_1525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1527 = i == 10'h2b ? _GEN_1526 : _GEN_1525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1528 = ~io_inputBit ? 1'h0 : _GEN_1527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1529 = i == 10'h30 ? _GEN_1528 : _GEN_1527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1530 = ~io_inputBit ? 1'h0 : _GEN_1529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1531 = i == 10'h58 ? _GEN_1530 : _GEN_1529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1532 = io_inputBit | _GEN_1531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1533 = i == 10'h58 ? _GEN_1532 : _GEN_1531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1534 = ~io_inputBit ? 1'h0 : _GEN_1533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1535 = i == 10'h59 ? _GEN_1534 : _GEN_1533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1536 = io_inputBit | _GEN_1535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1537 = i == 10'h59 ? _GEN_1536 : _GEN_1535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1538 = ~io_inputBit ? 1'h0 : _GEN_1537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1539 = i == 10'h5a ? _GEN_1538 : _GEN_1537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1540 = io_inputBit | _GEN_1539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1541 = i == 10'h5a ? _GEN_1540 : _GEN_1539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1542 = ~io_inputBit ? 1'h0 : _GEN_1541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1543 = i == 10'h5b ? _GEN_1542 : _GEN_1541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1544 = io_inputBit | _GEN_1543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1545 = i == 10'h5b ? _GEN_1544 : _GEN_1543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1546 = ~io_inputBit ? 1'h0 : _GEN_1545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1547 = i == 10'h5c ? _GEN_1546 : _GEN_1545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1548 = io_inputBit | _GEN_1547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1549 = i == 10'h5c ? _GEN_1548 : _GEN_1547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1550 = ~io_inputBit ? 1'h0 : _GEN_1549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1551 = i == 10'hc5 ? _GEN_1550 : _GEN_1549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1552 = io_inputBit | _GEN_1551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1553 = i == 10'hc5 ? _GEN_1552 : _GEN_1551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1554 = ~io_inputBit | _GEN_1553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1555 = i == 10'hc6 ? _GEN_1554 : _GEN_1553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1556 = io_inputBit ? 1'h0 : _GEN_1555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1557 = i == 10'hc6 ? _GEN_1556 : _GEN_1555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1558 = ~io_inputBit ? 1'h0 : _GEN_1557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1559 = i == 10'hc7 ? _GEN_1558 : _GEN_1557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1560 = io_inputBit | _GEN_1559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1561 = i == 10'hc7 ? _GEN_1560 : _GEN_1559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1562 = ~io_inputBit | _GEN_1561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1563 = i == 10'hc8 ? _GEN_1562 : _GEN_1561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1564 = io_inputBit ? 1'h0 : _GEN_1563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1565 = i == 10'hc8 ? _GEN_1564 : _GEN_1563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1566 = ~io_inputBit ? 1'h0 : _GEN_1565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1567 = i == 10'hc9 ? _GEN_1566 : _GEN_1565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1568 = io_inputBit | _GEN_1567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1569 = i == 10'hc9 ? _GEN_1568 : _GEN_1567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1570 = ~io_inputBit | _GEN_1569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1571 = i == 10'hca ? _GEN_1570 : _GEN_1569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1572 = io_inputBit ? 1'h0 : _GEN_1571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1573 = i == 10'hca ? _GEN_1572 : _GEN_1571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1574 = ~io_inputBit ? 1'h0 : _GEN_1573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1575 = i == 10'hcb ? _GEN_1574 : _GEN_1573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1576 = io_inputBit | _GEN_1575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1577 = i == 10'hcb ? _GEN_1576 : _GEN_1575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1578 = ~io_inputBit | _GEN_1577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1579 = i == 10'hcc ? _GEN_1578 : _GEN_1577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1580 = io_inputBit ? 1'h0 : _GEN_1579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1581 = i == 10'hcc ? _GEN_1580 : _GEN_1579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1582 = ~io_inputBit ? 1'h0 : _GEN_1581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1583 = i == 10'hcd ? _GEN_1582 : _GEN_1581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1584 = io_inputBit | _GEN_1583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1585 = i == 10'hcd ? _GEN_1584 : _GEN_1583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1586 = ~io_inputBit | _GEN_1585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1587 = i == 10'hce ? _GEN_1586 : _GEN_1585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1588 = io_inputBit ? 1'h0 : _GEN_1587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1589 = i == 10'hce ? _GEN_1588 : _GEN_1587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1590 = ~io_inputBit ? 1'h0 : _GEN_1209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1591 = i == 10'h1 ? _GEN_1590 : _GEN_1209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1592 = io_inputBit ? 1'h0 : _GEN_1591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1593 = i == 10'h2 ? _GEN_1592 : _GEN_1591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1594 = ~io_inputBit ? 1'h0 : _GEN_1593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1595 = i == 10'h4 ? _GEN_1594 : _GEN_1593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1596 = io_inputBit ? 1'h0 : _GEN_1595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1597 = i == 10'h5 ? _GEN_1596 : _GEN_1595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1598 = io_inputBit ? 1'h0 : _GEN_1597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1599 = i == 10'h16 ? _GEN_1598 : _GEN_1597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1600 = ~io_inputBit ? 1'h0 : _GEN_1599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1601 = i == 10'h17 ? _GEN_1600 : _GEN_1599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1602 = ~io_inputBit ? 1'h0 : _GEN_1601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1603 = i == 10'h2b ? _GEN_1602 : _GEN_1601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1604 = ~io_inputBit ? 1'h0 : _GEN_1603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1605 = i == 10'h30 ? _GEN_1604 : _GEN_1603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1606 = ~io_inputBit ? 1'h0 : _GEN_1605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1607 = i == 10'hb1 ? _GEN_1606 : _GEN_1605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1608 = io_inputBit | _GEN_1607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1609 = i == 10'hb1 ? _GEN_1608 : _GEN_1607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1610 = ~io_inputBit ? 1'h0 : _GEN_1609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1611 = i == 10'hb2 ? _GEN_1610 : _GEN_1609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1612 = io_inputBit | _GEN_1611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1613 = i == 10'hb2 ? _GEN_1612 : _GEN_1611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1614 = ~io_inputBit ? 1'h0 : _GEN_1613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1615 = i == 10'hb3 ? _GEN_1614 : _GEN_1613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1616 = io_inputBit | _GEN_1615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1617 = i == 10'hb3 ? _GEN_1616 : _GEN_1615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1618 = ~io_inputBit ? 1'h0 : _GEN_1617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1619 = i == 10'hb4 ? _GEN_1618 : _GEN_1617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1620 = io_inputBit | _GEN_1619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1621 = i == 10'hb4 ? _GEN_1620 : _GEN_1619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1622 = ~io_inputBit ? 1'h0 : _GEN_1621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1623 = i == 10'hb5 ? _GEN_1622 : _GEN_1621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1624 = io_inputBit | _GEN_1623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1625 = i == 10'hb5 ? _GEN_1624 : _GEN_1623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1626 = ~io_inputBit ? 1'h0 : _GEN_1625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1627 = i == 10'hb6 ? _GEN_1626 : _GEN_1625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1628 = io_inputBit | _GEN_1627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1629 = i == 10'hb6 ? _GEN_1628 : _GEN_1627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1630 = ~io_inputBit ? 1'h0 : _GEN_1629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1631 = i == 10'hb7 ? _GEN_1630 : _GEN_1629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1632 = io_inputBit | _GEN_1631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1633 = i == 10'hb7 ? _GEN_1632 : _GEN_1631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1634 = ~io_inputBit ? 1'h0 : _GEN_1633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1635 = i == 10'hb8 ? _GEN_1634 : _GEN_1633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1636 = io_inputBit | _GEN_1635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1637 = i == 10'hb8 ? _GEN_1636 : _GEN_1635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1638 = ~io_inputBit ? 1'h0 : _GEN_1637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1639 = i == 10'hb9 ? _GEN_1638 : _GEN_1637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1640 = io_inputBit | _GEN_1639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1641 = i == 10'hb9 ? _GEN_1640 : _GEN_1639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1642 = ~io_inputBit ? 1'h0 : _GEN_1641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1643 = i == 10'hba ? _GEN_1642 : _GEN_1641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1644 = io_inputBit | _GEN_1643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1645 = i == 10'hba ? _GEN_1644 : _GEN_1643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1646 = ~io_inputBit ? 1'h0 : _GEN_1645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1647 = i == 10'hc5 ? _GEN_1646 : _GEN_1645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1648 = io_inputBit | _GEN_1647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1649 = i == 10'hc5 ? _GEN_1648 : _GEN_1647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1650 = ~io_inputBit ? 1'h0 : _GEN_1649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1651 = i == 10'hc6 ? _GEN_1650 : _GEN_1649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1652 = io_inputBit | _GEN_1651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1653 = i == 10'hc6 ? _GEN_1652 : _GEN_1651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1654 = ~io_inputBit ? 1'h0 : _GEN_1653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1655 = i == 10'hc7 ? _GEN_1654 : _GEN_1653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1656 = io_inputBit | _GEN_1655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1657 = i == 10'hc7 ? _GEN_1656 : _GEN_1655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1658 = ~io_inputBit ? 1'h0 : _GEN_1657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1659 = i == 10'hc8 ? _GEN_1658 : _GEN_1657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1660 = io_inputBit | _GEN_1659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1661 = i == 10'hc8 ? _GEN_1660 : _GEN_1659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1662 = ~io_inputBit ? 1'h0 : _GEN_1661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1663 = i == 10'hc9 ? _GEN_1662 : _GEN_1661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1664 = io_inputBit | _GEN_1663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1665 = i == 10'hc9 ? _GEN_1664 : _GEN_1663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1666 = ~io_inputBit ? 1'h0 : _GEN_1665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1667 = i == 10'hca ? _GEN_1666 : _GEN_1665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1668 = io_inputBit | _GEN_1667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1669 = i == 10'hca ? _GEN_1668 : _GEN_1667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1670 = ~io_inputBit ? 1'h0 : _GEN_1669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1671 = i == 10'hcb ? _GEN_1670 : _GEN_1669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1672 = io_inputBit | _GEN_1671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1673 = i == 10'hcb ? _GEN_1672 : _GEN_1671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1674 = ~io_inputBit ? 1'h0 : _GEN_1673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1675 = i == 10'hcc ? _GEN_1674 : _GEN_1673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1676 = io_inputBit | _GEN_1675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1677 = i == 10'hcc ? _GEN_1676 : _GEN_1675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1678 = ~io_inputBit ? 1'h0 : _GEN_1677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1679 = i == 10'hcd ? _GEN_1678 : _GEN_1677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1680 = io_inputBit | _GEN_1679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1681 = i == 10'hcd ? _GEN_1680 : _GEN_1679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1682 = ~io_inputBit ? 1'h0 : _GEN_1681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1683 = i == 10'hce ? _GEN_1682 : _GEN_1681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1684 = io_inputBit | _GEN_1683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1685 = i == 10'hce ? _GEN_1684 : _GEN_1683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1686 = ~io_inputBit ? 1'h0 : _GEN_1237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1687 = i == 10'h0 ? _GEN_1686 : _GEN_1237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1688 = io_inputBit | _GEN_1687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1689 = i == 10'h2 ? _GEN_1688 : _GEN_1687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1690 = io_inputBit | _GEN_1689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1691 = i == 10'h5 ? _GEN_1690 : _GEN_1689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1692 = ~io_inputBit ? 1'h0 : _GEN_1691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1693 = i == 10'hb ? _GEN_1692 : _GEN_1691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1694 = ~io_inputBit ? 1'h0 : _GEN_1693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1695 = i == 10'h18 ? _GEN_1694 : _GEN_1693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1696 = io_inputBit | _GEN_1695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1697 = i == 10'h32 ? _GEN_1696 : _GEN_1695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1698 = io_inputBit | _GEN_1697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1699 = i == 10'h65 ? _GEN_1698 : _GEN_1697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1700 = ~io_inputBit ? 1'h0 : _GEN_1699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1701 = i == 10'hcb ? _GEN_1700 : _GEN_1699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1702 = io_inputBit | _GEN_1701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1703 = i == 10'hcb ? _GEN_1702 : _GEN_1701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1704 = ~io_inputBit ? 1'h0 : _GEN_1285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1705 = i == 10'h0 ? _GEN_1704 : _GEN_1285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1706 = io_inputBit | _GEN_1705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1707 = i == 10'h2 ? _GEN_1706 : _GEN_1705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1708 = io_inputBit | _GEN_1707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1709 = i == 10'h5 ? _GEN_1708 : _GEN_1707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1710 = ~io_inputBit ? 1'h0 : _GEN_1709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1711 = i == 10'hb ? _GEN_1710 : _GEN_1709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1712 = io_inputBit | _GEN_1711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1713 = i == 10'h31 ? _GEN_1712 : _GEN_1711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1714 = io_inputBit ? 1'h0 : _GEN_1713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1715 = i == 10'h32 ? _GEN_1714 : _GEN_1713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1716 = ~io_inputBit ? 1'h0 : _GEN_1715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1717 = i == 10'h63 ? _GEN_1716 : _GEN_1715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1718 = io_inputBit ? 1'h0 : _GEN_1717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1719 = i == 10'h65 ? _GEN_1718 : _GEN_1717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1720 = ~io_inputBit ? 1'h0 : _GEN_1719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1721 = i == 10'hc8 ? _GEN_1720 : _GEN_1719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1722 = io_inputBit | _GEN_1721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1723 = i == 10'hc8 ? _GEN_1722 : _GEN_1721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1724 = ~io_inputBit | _GEN_1723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1725 = i == 10'hcb ? _GEN_1724 : _GEN_1723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1726 = io_inputBit ? 1'h0 : _GEN_1725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1727 = i == 10'hcb ? _GEN_1726 : _GEN_1725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1728 = ~io_inputBit ? 1'h0 : _GEN_1347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1729 = i == 10'h0 ? _GEN_1728 : _GEN_1347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1730 = io_inputBit ? 1'h0 : _GEN_1729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1731 = i == 10'h2 ? _GEN_1730 : _GEN_1729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1732 = io_inputBit ? 1'h0 : _GEN_1731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1733 = i == 10'h5 ? _GEN_1732 : _GEN_1731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1734 = ~io_inputBit ? 1'h0 : _GEN_1733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1735 = i == 10'hb ? _GEN_1734 : _GEN_1733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1736 = io_inputBit | _GEN_1735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1737 = i == 10'h32 ? _GEN_1736 : _GEN_1735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1738 = ~io_inputBit | _GEN_1737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1739 = i == 10'h63 ? _GEN_1738 : _GEN_1737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1740 = ~io_inputBit ? 1'h0 : _GEN_1739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1741 = i == 10'h64 ? _GEN_1740 : _GEN_1739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1742 = io_inputBit | _GEN_1741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1743 = i == 10'h64 ? _GEN_1742 : _GEN_1741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1744 = io_inputBit ? 1'h0 : _GEN_1743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1745 = i == 10'h65 ? _GEN_1744 : _GEN_1743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1746 = ~io_inputBit | _GEN_1745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1747 = i == 10'hc8 ? _GEN_1746 : _GEN_1745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1748 = io_inputBit ? 1'h0 : _GEN_1747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1749 = i == 10'hc8 ? _GEN_1748 : _GEN_1747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1750 = ~io_inputBit | _GEN_1749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1751 = i == 10'hcb ? _GEN_1750 : _GEN_1749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1752 = io_inputBit ? 1'h0 : _GEN_1751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1753 = i == 10'hcb ? _GEN_1752 : _GEN_1751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1754 = ~io_inputBit ? 1'h0 : _GEN_1427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1755 = i == 10'h0 ? _GEN_1754 : _GEN_1427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1756 = io_inputBit ? 1'h0 : _GEN_1755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1757 = i == 10'h2 ? _GEN_1756 : _GEN_1755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1758 = io_inputBit ? 1'h0 : _GEN_1757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1759 = i == 10'h5 ? _GEN_1758 : _GEN_1757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1760 = ~io_inputBit ? 1'h0 : _GEN_1759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1761 = i == 10'h17 ? _GEN_1760 : _GEN_1759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1762 = ~io_inputBit ? 1'h0 : _GEN_1761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1763 = i == 10'h30 ? _GEN_1762 : _GEN_1761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1764 = ~io_inputBit ? 1'h0 : _GEN_1763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1765 = i == 10'h62 ? _GEN_1764 : _GEN_1763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1766 = io_inputBit | _GEN_1765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1767 = i == 10'h62 ? _GEN_1766 : _GEN_1765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1768 = ~io_inputBit | _GEN_1767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1769 = i == 10'h64 ? _GEN_1768 : _GEN_1767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1770 = io_inputBit ? 1'h0 : _GEN_1769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1771 = i == 10'h64 ? _GEN_1770 : _GEN_1769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1772 = ~io_inputBit ? 1'h0 : _GEN_1771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1773 = i == 10'h66 ? _GEN_1772 : _GEN_1771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1774 = io_inputBit | _GEN_1773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1775 = i == 10'h66 ? _GEN_1774 : _GEN_1773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1776 = ~io_inputBit ? 1'h0 : _GEN_1775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1777 = i == 10'hc7 ? _GEN_1776 : _GEN_1775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1778 = io_inputBit | _GEN_1777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1779 = i == 10'hc7 ? _GEN_1778 : _GEN_1777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1780 = ~io_inputBit | _GEN_1779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1781 = i == 10'hc8 ? _GEN_1780 : _GEN_1779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1782 = io_inputBit ? 1'h0 : _GEN_1781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1783 = i == 10'hc8 ? _GEN_1782 : _GEN_1781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1784 = ~io_inputBit | _GEN_1783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1785 = i == 10'hcb ? _GEN_1784 : _GEN_1783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1786 = io_inputBit ? 1'h0 : _GEN_1785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1787 = i == 10'hcb ? _GEN_1786 : _GEN_1785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1788 = ~io_inputBit ? 1'h0 : _GEN_1787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1789 = i == 10'hcc ? _GEN_1788 : _GEN_1787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1790 = io_inputBit | _GEN_1789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1791 = i == 10'hcc ? _GEN_1790 : _GEN_1789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1792 = ~io_inputBit ? 1'h0 : _GEN_1513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1793 = i == 10'h0 ? _GEN_1792 : _GEN_1513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1794 = io_inputBit | _GEN_1793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1795 = i == 10'h2 ? _GEN_1794 : _GEN_1793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1796 = io_inputBit | _GEN_1795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1797 = i == 10'h5 ? _GEN_1796 : _GEN_1795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1798 = ~io_inputBit ? 1'h0 : _GEN_1797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1799 = i == 10'h17 ? _GEN_1798 : _GEN_1797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1800 = ~io_inputBit ? 1'h0 : _GEN_1799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1801 = i == 10'h30 ? _GEN_1800 : _GEN_1799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1802 = ~io_inputBit ? 1'h0 : _GEN_1801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1803 = i == 10'hc5 ? _GEN_1802 : _GEN_1801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1804 = io_inputBit | _GEN_1803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1805 = i == 10'hc5 ? _GEN_1804 : _GEN_1803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1806 = ~io_inputBit ? 1'h0 : _GEN_1805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1807 = i == 10'hc6 ? _GEN_1806 : _GEN_1805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1808 = io_inputBit | _GEN_1807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1809 = i == 10'hc6 ? _GEN_1808 : _GEN_1807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1810 = ~io_inputBit | _GEN_1809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1811 = i == 10'hc7 ? _GEN_1810 : _GEN_1809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1812 = io_inputBit ? 1'h0 : _GEN_1811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1813 = i == 10'hc7 ? _GEN_1812 : _GEN_1811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1814 = ~io_inputBit | _GEN_1813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1815 = i == 10'hc8 ? _GEN_1814 : _GEN_1813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1816 = io_inputBit ? 1'h0 : _GEN_1815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1817 = i == 10'hc8 ? _GEN_1816 : _GEN_1815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1818 = ~io_inputBit ? 1'h0 : _GEN_1817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1819 = i == 10'hc9 ? _GEN_1818 : _GEN_1817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1820 = io_inputBit | _GEN_1819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1821 = i == 10'hc9 ? _GEN_1820 : _GEN_1819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1822 = ~io_inputBit ? 1'h0 : _GEN_1821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1823 = i == 10'hca ? _GEN_1822 : _GEN_1821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1824 = io_inputBit | _GEN_1823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1825 = i == 10'hca ? _GEN_1824 : _GEN_1823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1826 = ~io_inputBit | _GEN_1825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1827 = i == 10'hcb ? _GEN_1826 : _GEN_1825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1828 = io_inputBit ? 1'h0 : _GEN_1827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1829 = i == 10'hcb ? _GEN_1828 : _GEN_1827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1830 = ~io_inputBit | _GEN_1829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1831 = i == 10'hcc ? _GEN_1830 : _GEN_1829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1832 = io_inputBit ? 1'h0 : _GEN_1831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1833 = i == 10'hcc ? _GEN_1832 : _GEN_1831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1834 = ~io_inputBit ? 1'h0 : _GEN_1833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1835 = i == 10'hcd ? _GEN_1834 : _GEN_1833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1836 = io_inputBit | _GEN_1835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1837 = i == 10'hcd ? _GEN_1836 : _GEN_1835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1838 = ~io_inputBit ? 1'h0 : _GEN_1837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1839 = i == 10'hce ? _GEN_1838 : _GEN_1837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1840 = io_inputBit | _GEN_1839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1841 = i == 10'hce ? _GEN_1840 : _GEN_1839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1842 = ~io_inputBit ? 1'h0 : _GEN_1589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1843 = i == 10'h0 ? _GEN_1842 : _GEN_1589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1844 = io_inputBit ? 1'h0 : _GEN_1843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1845 = i == 10'h2 ? _GEN_1844 : _GEN_1843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1846 = io_inputBit ? 1'h0 : _GEN_1845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1847 = i == 10'h5 ? _GEN_1846 : _GEN_1845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1848 = ~io_inputBit ? 1'h0 : _GEN_1847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1849 = i == 10'h17 ? _GEN_1848 : _GEN_1847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1850 = ~io_inputBit ? 1'h0 : _GEN_1849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1851 = i == 10'h30 ? _GEN_1850 : _GEN_1849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1852 = ~io_inputBit ? 1'h0 : _GEN_1851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1853 = i == 10'h62 ? _GEN_1852 : _GEN_1851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1854 = io_inputBit | _GEN_1853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1855 = i == 10'h62 ? _GEN_1854 : _GEN_1853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1856 = ~io_inputBit ? 1'h0 : _GEN_1855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1857 = i == 10'h63 ? _GEN_1856 : _GEN_1855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1858 = io_inputBit | _GEN_1857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1859 = i == 10'h63 ? _GEN_1858 : _GEN_1857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1860 = ~io_inputBit ? 1'h0 : _GEN_1859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1861 = i == 10'h64 ? _GEN_1860 : _GEN_1859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1862 = io_inputBit | _GEN_1861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1863 = i == 10'h64 ? _GEN_1862 : _GEN_1861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1864 = ~io_inputBit ? 1'h0 : _GEN_1863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1865 = i == 10'h65 ? _GEN_1864 : _GEN_1863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1866 = io_inputBit | _GEN_1865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1867 = i == 10'h65 ? _GEN_1866 : _GEN_1865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1868 = ~io_inputBit ? 1'h0 : _GEN_1867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1869 = i == 10'h66 ? _GEN_1868 : _GEN_1867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1870 = io_inputBit | _GEN_1869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1871 = i == 10'h66 ? _GEN_1870 : _GEN_1869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1872 = ~io_inputBit ? 1'h0 : _GEN_1685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1873 = i == 10'h0 ? _GEN_1872 : _GEN_1685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1874 = io_inputBit ? 1'h0 : _GEN_1873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1875 = i == 10'h2 ? _GEN_1874 : _GEN_1873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1876 = io_inputBit ? 1'h0 : _GEN_1875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1877 = i == 10'h5 ? _GEN_1876 : _GEN_1875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1878 = ~io_inputBit ? 1'h0 : _GEN_1877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1879 = i == 10'h17 ? _GEN_1878 : _GEN_1877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1880 = ~io_inputBit ? 1'h0 : _GEN_1879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1881 = i == 10'h30 ? _GEN_1880 : _GEN_1879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1882 = ~io_inputBit ? 1'h0 : _GEN_1881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1883 = i == 10'hc5 ? _GEN_1882 : _GEN_1881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1884 = io_inputBit | _GEN_1883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1885 = i == 10'hc5 ? _GEN_1884 : _GEN_1883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1886 = ~io_inputBit ? 1'h0 : _GEN_1885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1887 = i == 10'hc6 ? _GEN_1886 : _GEN_1885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1888 = io_inputBit | _GEN_1887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1889 = i == 10'hc6 ? _GEN_1888 : _GEN_1887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1890 = ~io_inputBit ? 1'h0 : _GEN_1889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1891 = i == 10'hc7 ? _GEN_1890 : _GEN_1889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1892 = io_inputBit | _GEN_1891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1893 = i == 10'hc7 ? _GEN_1892 : _GEN_1891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1894 = ~io_inputBit ? 1'h0 : _GEN_1893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1895 = i == 10'hc8 ? _GEN_1894 : _GEN_1893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1896 = io_inputBit | _GEN_1895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1897 = i == 10'hc8 ? _GEN_1896 : _GEN_1895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1898 = ~io_inputBit ? 1'h0 : _GEN_1897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1899 = i == 10'hc9 ? _GEN_1898 : _GEN_1897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1900 = io_inputBit | _GEN_1899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1901 = i == 10'hc9 ? _GEN_1900 : _GEN_1899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1902 = ~io_inputBit ? 1'h0 : _GEN_1901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1903 = i == 10'hca ? _GEN_1902 : _GEN_1901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1904 = io_inputBit | _GEN_1903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1905 = i == 10'hca ? _GEN_1904 : _GEN_1903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1906 = ~io_inputBit ? 1'h0 : _GEN_1905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1907 = i == 10'hcb ? _GEN_1906 : _GEN_1905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1908 = io_inputBit | _GEN_1907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1909 = i == 10'hcb ? _GEN_1908 : _GEN_1907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1910 = ~io_inputBit ? 1'h0 : _GEN_1909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1911 = i == 10'hcc ? _GEN_1910 : _GEN_1909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1912 = io_inputBit | _GEN_1911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1913 = i == 10'hcc ? _GEN_1912 : _GEN_1911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1914 = ~io_inputBit ? 1'h0 : _GEN_1913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1915 = i == 10'hcd ? _GEN_1914 : _GEN_1913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1916 = io_inputBit | _GEN_1915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1917 = i == 10'hcd ? _GEN_1916 : _GEN_1915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1918 = ~io_inputBit ? 1'h0 : _GEN_1917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1919 = i == 10'hce ? _GEN_1918 : _GEN_1917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1920 = io_inputBit | _GEN_1919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1921 = i == 10'hce ? _GEN_1920 : _GEN_1919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1922 = io_inputBit ? 1'h0 : _GEN_1703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1923 = i == 10'h0 ? _GEN_1922 : _GEN_1703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1924 = io_inputBit ? 1'h0 : _GEN_1923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1925 = i == 10'h1 ? _GEN_1924 : _GEN_1923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1926 = io_inputBit ? 1'h0 : _GEN_1925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1927 = i == 10'h3 ? _GEN_1926 : _GEN_1925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1928 = ~io_inputBit | _GEN_1927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1929 = i == 10'h7 ? _GEN_1928 : _GEN_1927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1930 = io_inputBit ? 1'h0 : _GEN_1929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1931 = i == 10'h10 ? _GEN_1930 : _GEN_1929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1932 = ~io_inputBit | _GEN_1931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1933 = i == 10'h21 ? _GEN_1932 : _GEN_1931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1934 = io_inputBit ? 1'h0 : _GEN_1933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1935 = i == 10'h44 ? _GEN_1934 : _GEN_1933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1936 = ~io_inputBit | _GEN_1935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1937 = i == 10'h89 ? _GEN_1936 : _GEN_1935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1938 = ~io_inputBit | _GEN_1937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1939 = i == 10'h114 ? _GEN_1938 : _GEN_1937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1940 = ~io_inputBit | _GEN_1939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1941 = i == 10'h22a ? _GEN_1940 : _GEN_1939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1942 = io_inputBit ? 1'h0 : _GEN_1941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1943 = i == 10'h22a ? _GEN_1942 : _GEN_1941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1944 = io_inputBit ? 1'h0 : _GEN_1727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1945 = i == 10'h0 ? _GEN_1944 : _GEN_1727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1946 = io_inputBit ? 1'h0 : _GEN_1945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1947 = i == 10'h1 ? _GEN_1946 : _GEN_1945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1948 = io_inputBit ? 1'h0 : _GEN_1947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1949 = i == 10'h3 ? _GEN_1948 : _GEN_1947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1950 = ~io_inputBit | _GEN_1949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1951 = i == 10'hf ? _GEN_1950 : _GEN_1949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1952 = ~io_inputBit | _GEN_1951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1953 = i == 10'h20 ? _GEN_1952 : _GEN_1951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1954 = ~io_inputBit ? 1'h0 : _GEN_1953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1955 = i == 10'h21 ? _GEN_1954 : _GEN_1953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1956 = ~io_inputBit | _GEN_1955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1957 = i == 10'h22 ? _GEN_1956 : _GEN_1955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1958 = io_inputBit ? 1'h0 : _GEN_1957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1959 = i == 10'h42 ? _GEN_1958 : _GEN_1957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1960 = io_inputBit | _GEN_1959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1961 = i == 10'h44 ? _GEN_1960 : _GEN_1959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1962 = io_inputBit ? 1'h0 : _GEN_1961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1963 = i == 10'h46 ? _GEN_1962 : _GEN_1961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1964 = ~io_inputBit | _GEN_1963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1965 = i == 10'h85 ? _GEN_1964 : _GEN_1963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1966 = ~io_inputBit ? 1'h0 : _GEN_1965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1967 = i == 10'h89 ? _GEN_1966 : _GEN_1965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1968 = ~io_inputBit | _GEN_1967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1969 = i == 10'h8d ? _GEN_1968 : _GEN_1967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1970 = ~io_inputBit | _GEN_1969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1971 = i == 10'h10c ? _GEN_1970 : _GEN_1969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1972 = ~io_inputBit ? 1'h0 : _GEN_1971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1973 = i == 10'h114 ? _GEN_1972 : _GEN_1971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1974 = ~io_inputBit | _GEN_1973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1975 = i == 10'h11c ? _GEN_1974 : _GEN_1973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1976 = ~io_inputBit | _GEN_1975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1977 = i == 10'h21a ? _GEN_1976 : _GEN_1975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1978 = io_inputBit ? 1'h0 : _GEN_1977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1979 = i == 10'h21a ? _GEN_1978 : _GEN_1977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1980 = ~io_inputBit ? 1'h0 : _GEN_1979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1981 = i == 10'h22a ? _GEN_1980 : _GEN_1979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1982 = io_inputBit | _GEN_1981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1983 = i == 10'h22a ? _GEN_1982 : _GEN_1981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1984 = ~io_inputBit | _GEN_1983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1985 = i == 10'h23a ? _GEN_1984 : _GEN_1983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1986 = io_inputBit ? 1'h0 : _GEN_1985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1987 = i == 10'h23a ? _GEN_1986 : _GEN_1985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1988 = io_inputBit ? 1'h0 : _GEN_1753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1989 = i == 10'h0 ? _GEN_1988 : _GEN_1753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1990 = io_inputBit ? 1'h0 : _GEN_1989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1991 = i == 10'h1 ? _GEN_1990 : _GEN_1989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1992 = io_inputBit ? 1'h0 : _GEN_1991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1993 = i == 10'h8 ? _GEN_1992 : _GEN_1991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1994 = ~io_inputBit ? 1'h0 : _GEN_1993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1995 = i == 10'hf ? _GEN_1994 : _GEN_1993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1996 = io_inputBit ? 1'h0 : _GEN_1995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1997 = i == 10'h11 ? _GEN_1996 : _GEN_1995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1998 = ~io_inputBit ? 1'h0 : _GEN_1997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1999 = i == 10'h20 ? _GEN_1998 : _GEN_1997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2000 = io_inputBit ? 1'h0 : _GEN_1999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2001 = i == 10'h23 ? _GEN_2000 : _GEN_1999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2002 = io_inputBit | _GEN_2001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2003 = i == 10'h42 ? _GEN_2002 : _GEN_2001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2004 = io_inputBit ? 1'h0 : _GEN_2003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2005 = i == 10'h43 ? _GEN_2004 : _GEN_2003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2006 = io_inputBit | _GEN_2005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2007 = i == 10'h44 ? _GEN_2006 : _GEN_2005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2008 = io_inputBit ? 1'h0 : _GEN_2007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2009 = i == 10'h45 ? _GEN_2008 : _GEN_2007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2010 = io_inputBit | _GEN_2009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2011 = i == 10'h46 ? _GEN_2010 : _GEN_2009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2012 = io_inputBit ? 1'h0 : _GEN_2011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2013 = i == 10'h47 ? _GEN_2012 : _GEN_2011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2014 = ~io_inputBit ? 1'h0 : _GEN_2013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2015 = i == 10'h85 ? _GEN_2014 : _GEN_2013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2016 = ~io_inputBit | _GEN_2015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2017 = i == 10'h87 ? _GEN_2016 : _GEN_2015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2018 = ~io_inputBit ? 1'h0 : _GEN_2017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2019 = i == 10'h89 ? _GEN_2018 : _GEN_2017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2020 = ~io_inputBit | _GEN_2019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2021 = i == 10'h8b ? _GEN_2020 : _GEN_2019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2022 = ~io_inputBit ? 1'h0 : _GEN_2021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2023 = i == 10'h8d ? _GEN_2022 : _GEN_2021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2024 = ~io_inputBit | _GEN_2023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2025 = i == 10'h8f ? _GEN_2024 : _GEN_2023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2026 = ~io_inputBit ? 1'h0 : _GEN_2025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2027 = i == 10'h10c ? _GEN_2026 : _GEN_2025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2028 = ~io_inputBit | _GEN_2027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2029 = i == 10'h110 ? _GEN_2028 : _GEN_2027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2030 = ~io_inputBit ? 1'h0 : _GEN_2029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2031 = i == 10'h114 ? _GEN_2030 : _GEN_2029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2032 = ~io_inputBit | _GEN_2031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2033 = i == 10'h118 ? _GEN_2032 : _GEN_2031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2034 = ~io_inputBit ? 1'h0 : _GEN_2033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2035 = i == 10'h11c ? _GEN_2034 : _GEN_2033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2036 = ~io_inputBit | _GEN_2035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2037 = i == 10'h120 ? _GEN_2036 : _GEN_2035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2038 = ~io_inputBit ? 1'h0 : _GEN_2037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2039 = i == 10'h21a ? _GEN_2038 : _GEN_2037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2040 = io_inputBit | _GEN_2039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2041 = i == 10'h21a ? _GEN_2040 : _GEN_2039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2042 = ~io_inputBit | _GEN_2041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2043 = i == 10'h222 ? _GEN_2042 : _GEN_2041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2044 = io_inputBit ? 1'h0 : _GEN_2043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2045 = i == 10'h222 ? _GEN_2044 : _GEN_2043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2046 = ~io_inputBit ? 1'h0 : _GEN_2045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2047 = i == 10'h22a ? _GEN_2046 : _GEN_2045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2048 = io_inputBit | _GEN_2047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2049 = i == 10'h22a ? _GEN_2048 : _GEN_2047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2050 = ~io_inputBit | _GEN_2049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2051 = i == 10'h232 ? _GEN_2050 : _GEN_2049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2052 = io_inputBit ? 1'h0 : _GEN_2051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2053 = i == 10'h232 ? _GEN_2052 : _GEN_2051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2054 = ~io_inputBit ? 1'h0 : _GEN_2053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2055 = i == 10'h23a ? _GEN_2054 : _GEN_2053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2056 = io_inputBit | _GEN_2055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2057 = i == 10'h23a ? _GEN_2056 : _GEN_2055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2058 = ~io_inputBit | _GEN_2057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2059 = i == 10'h242 ? _GEN_2058 : _GEN_2057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2060 = io_inputBit ? 1'h0 : _GEN_2059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2061 = i == 10'h242 ? _GEN_2060 : _GEN_2059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2062 = io_inputBit ? 1'h0 : _GEN_1791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2063 = i == 10'h0 ? _GEN_2062 : _GEN_1791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2064 = io_inputBit ? 1'h0 : _GEN_2063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2065 = i == 10'h1 ? _GEN_2064 : _GEN_2063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2066 = io_inputBit ? 1'h0 : _GEN_2065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2067 = i == 10'h8 ? _GEN_2066 : _GEN_2065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2068 = ~io_inputBit ? 1'h0 : _GEN_2067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2069 = i == 10'hf ? _GEN_2068 : _GEN_2067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2070 = io_inputBit ? 1'h0 : _GEN_2069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2071 = i == 10'h11 ? _GEN_2070 : _GEN_2069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2072 = ~io_inputBit ? 1'h0 : _GEN_2071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2073 = i == 10'h20 ? _GEN_2072 : _GEN_2071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2074 = io_inputBit ? 1'h0 : _GEN_2073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2075 = i == 10'h23 ? _GEN_2074 : _GEN_2073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2076 = ~io_inputBit ? 1'h0 : _GEN_2075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2077 = i == 10'h85 ? _GEN_2076 : _GEN_2075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2078 = ~io_inputBit | _GEN_2077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2079 = i == 10'h86 ? _GEN_2078 : _GEN_2077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2080 = ~io_inputBit ? 1'h0 : _GEN_2079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2081 = i == 10'h87 ? _GEN_2080 : _GEN_2079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2082 = ~io_inputBit | _GEN_2081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2083 = i == 10'h88 ? _GEN_2082 : _GEN_2081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2084 = ~io_inputBit ? 1'h0 : _GEN_2083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2085 = i == 10'h89 ? _GEN_2084 : _GEN_2083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2086 = ~io_inputBit | _GEN_2085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2087 = i == 10'h8a ? _GEN_2086 : _GEN_2085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2088 = ~io_inputBit ? 1'h0 : _GEN_2087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2089 = i == 10'h8b ? _GEN_2088 : _GEN_2087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2090 = ~io_inputBit | _GEN_2089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2091 = i == 10'h8c ? _GEN_2090 : _GEN_2089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2092 = ~io_inputBit ? 1'h0 : _GEN_2091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2093 = i == 10'h8d ? _GEN_2092 : _GEN_2091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2094 = ~io_inputBit | _GEN_2093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2095 = i == 10'h8e ? _GEN_2094 : _GEN_2093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2096 = ~io_inputBit ? 1'h0 : _GEN_2095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2097 = i == 10'h8f ? _GEN_2096 : _GEN_2095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2098 = ~io_inputBit | _GEN_2097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2099 = i == 10'h90 ? _GEN_2098 : _GEN_2097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2100 = ~io_inputBit ? 1'h0 : _GEN_2099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2101 = i == 10'h10c ? _GEN_2100 : _GEN_2099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2102 = ~io_inputBit | _GEN_2101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2103 = i == 10'h10e ? _GEN_2102 : _GEN_2101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2104 = ~io_inputBit ? 1'h0 : _GEN_2103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2105 = i == 10'h110 ? _GEN_2104 : _GEN_2103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2106 = ~io_inputBit | _GEN_2105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2107 = i == 10'h112 ? _GEN_2106 : _GEN_2105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2108 = ~io_inputBit ? 1'h0 : _GEN_2107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2109 = i == 10'h114 ? _GEN_2108 : _GEN_2107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2110 = ~io_inputBit | _GEN_2109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2111 = i == 10'h116 ? _GEN_2110 : _GEN_2109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2112 = ~io_inputBit ? 1'h0 : _GEN_2111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2113 = i == 10'h118 ? _GEN_2112 : _GEN_2111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2114 = ~io_inputBit | _GEN_2113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2115 = i == 10'h11a ? _GEN_2114 : _GEN_2113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2116 = ~io_inputBit ? 1'h0 : _GEN_2115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2117 = i == 10'h11c ? _GEN_2116 : _GEN_2115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2118 = ~io_inputBit | _GEN_2117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2119 = i == 10'h11e ? _GEN_2118 : _GEN_2117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2120 = ~io_inputBit ? 1'h0 : _GEN_2119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2121 = i == 10'h120 ? _GEN_2120 : _GEN_2119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2122 = ~io_inputBit | _GEN_2121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2123 = i == 10'h122 ? _GEN_2122 : _GEN_2121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2124 = ~io_inputBit ? 1'h0 : _GEN_2123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2125 = i == 10'h21a ? _GEN_2124 : _GEN_2123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2126 = io_inputBit | _GEN_2125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2127 = i == 10'h21a ? _GEN_2126 : _GEN_2125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2128 = ~io_inputBit | _GEN_2127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2129 = i == 10'h21e ? _GEN_2128 : _GEN_2127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2130 = io_inputBit ? 1'h0 : _GEN_2129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2131 = i == 10'h21e ? _GEN_2130 : _GEN_2129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2132 = ~io_inputBit ? 1'h0 : _GEN_2131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2133 = i == 10'h222 ? _GEN_2132 : _GEN_2131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2134 = io_inputBit | _GEN_2133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2135 = i == 10'h222 ? _GEN_2134 : _GEN_2133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2136 = ~io_inputBit | _GEN_2135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2137 = i == 10'h226 ? _GEN_2136 : _GEN_2135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2138 = io_inputBit ? 1'h0 : _GEN_2137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2139 = i == 10'h226 ? _GEN_2138 : _GEN_2137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2140 = ~io_inputBit ? 1'h0 : _GEN_2139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2141 = i == 10'h22a ? _GEN_2140 : _GEN_2139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2142 = io_inputBit | _GEN_2141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2143 = i == 10'h22a ? _GEN_2142 : _GEN_2141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2144 = ~io_inputBit | _GEN_2143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2145 = i == 10'h22e ? _GEN_2144 : _GEN_2143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2146 = io_inputBit ? 1'h0 : _GEN_2145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2147 = i == 10'h22e ? _GEN_2146 : _GEN_2145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2148 = ~io_inputBit ? 1'h0 : _GEN_2147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2149 = i == 10'h232 ? _GEN_2148 : _GEN_2147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2150 = io_inputBit | _GEN_2149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2151 = i == 10'h232 ? _GEN_2150 : _GEN_2149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2152 = ~io_inputBit | _GEN_2151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2153 = i == 10'h236 ? _GEN_2152 : _GEN_2151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2154 = io_inputBit ? 1'h0 : _GEN_2153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2155 = i == 10'h236 ? _GEN_2154 : _GEN_2153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2156 = ~io_inputBit ? 1'h0 : _GEN_2155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2157 = i == 10'h23a ? _GEN_2156 : _GEN_2155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2158 = io_inputBit | _GEN_2157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2159 = i == 10'h23a ? _GEN_2158 : _GEN_2157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2160 = ~io_inputBit | _GEN_2159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2161 = i == 10'h23e ? _GEN_2160 : _GEN_2159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2162 = io_inputBit ? 1'h0 : _GEN_2161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2163 = i == 10'h23e ? _GEN_2162 : _GEN_2161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2164 = ~io_inputBit ? 1'h0 : _GEN_2163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2165 = i == 10'h242 ? _GEN_2164 : _GEN_2163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2166 = io_inputBit | _GEN_2165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2167 = i == 10'h242 ? _GEN_2166 : _GEN_2165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2168 = ~io_inputBit | _GEN_2167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2169 = i == 10'h246 ? _GEN_2168 : _GEN_2167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2170 = io_inputBit ? 1'h0 : _GEN_2169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2171 = i == 10'h246 ? _GEN_2170 : _GEN_2169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2172 = io_inputBit ? 1'h0 : _GEN_1841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2173 = i == 10'h0 ? _GEN_2172 : _GEN_1841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2174 = io_inputBit ? 1'h0 : _GEN_2173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2175 = i == 10'h1 ? _GEN_2174 : _GEN_2173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2176 = io_inputBit ? 1'h0 : _GEN_2175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2177 = i == 10'h8 ? _GEN_2176 : _GEN_2175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2178 = ~io_inputBit | _GEN_2177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2179 = i == 10'hf ? _GEN_2178 : _GEN_2177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2180 = io_inputBit ? 1'h0 : _GEN_2179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2181 = i == 10'h11 ? _GEN_2180 : _GEN_2179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2182 = ~io_inputBit | _GEN_2181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2183 = i == 10'h20 ? _GEN_2182 : _GEN_2181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2184 = io_inputBit ? 1'h0 : _GEN_2183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2185 = i == 10'h48 ? _GEN_2184 : _GEN_2183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2186 = io_inputBit ? 1'h0 : _GEN_2185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2187 = i == 10'h91 ? _GEN_2186 : _GEN_2185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2188 = ~io_inputBit | _GEN_2187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2189 = i == 10'h10b ? _GEN_2188 : _GEN_2187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2190 = ~io_inputBit ? 1'h0 : _GEN_2189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2191 = i == 10'h10c ? _GEN_2190 : _GEN_2189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2192 = ~io_inputBit | _GEN_2191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2193 = i == 10'h10d ? _GEN_2192 : _GEN_2191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2194 = ~io_inputBit ? 1'h0 : _GEN_2193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2195 = i == 10'h10e ? _GEN_2194 : _GEN_2193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2196 = ~io_inputBit | _GEN_2195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2197 = i == 10'h10f ? _GEN_2196 : _GEN_2195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2198 = ~io_inputBit ? 1'h0 : _GEN_2197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2199 = i == 10'h110 ? _GEN_2198 : _GEN_2197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2200 = ~io_inputBit | _GEN_2199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2201 = i == 10'h111 ? _GEN_2200 : _GEN_2199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2202 = ~io_inputBit ? 1'h0 : _GEN_2201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2203 = i == 10'h112 ? _GEN_2202 : _GEN_2201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2204 = ~io_inputBit | _GEN_2203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2205 = i == 10'h113 ? _GEN_2204 : _GEN_2203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2206 = ~io_inputBit ? 1'h0 : _GEN_2205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2207 = i == 10'h114 ? _GEN_2206 : _GEN_2205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2208 = ~io_inputBit | _GEN_2207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2209 = i == 10'h115 ? _GEN_2208 : _GEN_2207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2210 = ~io_inputBit ? 1'h0 : _GEN_2209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2211 = i == 10'h116 ? _GEN_2210 : _GEN_2209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2212 = ~io_inputBit | _GEN_2211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2213 = i == 10'h117 ? _GEN_2212 : _GEN_2211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2214 = ~io_inputBit ? 1'h0 : _GEN_2213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2215 = i == 10'h118 ? _GEN_2214 : _GEN_2213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2216 = ~io_inputBit | _GEN_2215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2217 = i == 10'h119 ? _GEN_2216 : _GEN_2215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2218 = ~io_inputBit ? 1'h0 : _GEN_2217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2219 = i == 10'h11a ? _GEN_2218 : _GEN_2217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2220 = ~io_inputBit | _GEN_2219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2221 = i == 10'h11b ? _GEN_2220 : _GEN_2219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2222 = ~io_inputBit ? 1'h0 : _GEN_2221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2223 = i == 10'h11c ? _GEN_2222 : _GEN_2221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2224 = ~io_inputBit | _GEN_2223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2225 = i == 10'h11d ? _GEN_2224 : _GEN_2223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2226 = ~io_inputBit ? 1'h0 : _GEN_2225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2227 = i == 10'h11e ? _GEN_2226 : _GEN_2225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2228 = ~io_inputBit | _GEN_2227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2229 = i == 10'h11f ? _GEN_2228 : _GEN_2227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2230 = ~io_inputBit ? 1'h0 : _GEN_2229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2231 = i == 10'h120 ? _GEN_2230 : _GEN_2229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2232 = ~io_inputBit | _GEN_2231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2233 = i == 10'h121 ? _GEN_2232 : _GEN_2231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2234 = ~io_inputBit ? 1'h0 : _GEN_2233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2235 = i == 10'h122 ? _GEN_2234 : _GEN_2233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2236 = ~io_inputBit | _GEN_2235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2237 = i == 10'h123 ? _GEN_2236 : _GEN_2235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2238 = ~io_inputBit | _GEN_2237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2239 = i == 10'h218 ? _GEN_2238 : _GEN_2237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2240 = io_inputBit ? 1'h0 : _GEN_2239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2241 = i == 10'h218 ? _GEN_2240 : _GEN_2239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2242 = ~io_inputBit ? 1'h0 : _GEN_2241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2243 = i == 10'h21a ? _GEN_2242 : _GEN_2241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2244 = io_inputBit | _GEN_2243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2245 = i == 10'h21a ? _GEN_2244 : _GEN_2243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2246 = ~io_inputBit | _GEN_2245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2247 = i == 10'h21c ? _GEN_2246 : _GEN_2245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2248 = io_inputBit ? 1'h0 : _GEN_2247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2249 = i == 10'h21c ? _GEN_2248 : _GEN_2247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2250 = ~io_inputBit ? 1'h0 : _GEN_2249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2251 = i == 10'h21e ? _GEN_2250 : _GEN_2249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2252 = io_inputBit | _GEN_2251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2253 = i == 10'h21e ? _GEN_2252 : _GEN_2251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2254 = ~io_inputBit | _GEN_2253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2255 = i == 10'h220 ? _GEN_2254 : _GEN_2253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2256 = io_inputBit ? 1'h0 : _GEN_2255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2257 = i == 10'h220 ? _GEN_2256 : _GEN_2255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2258 = ~io_inputBit ? 1'h0 : _GEN_2257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2259 = i == 10'h222 ? _GEN_2258 : _GEN_2257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2260 = io_inputBit | _GEN_2259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2261 = i == 10'h222 ? _GEN_2260 : _GEN_2259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2262 = ~io_inputBit | _GEN_2261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2263 = i == 10'h224 ? _GEN_2262 : _GEN_2261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2264 = io_inputBit ? 1'h0 : _GEN_2263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2265 = i == 10'h224 ? _GEN_2264 : _GEN_2263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2266 = ~io_inputBit ? 1'h0 : _GEN_2265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2267 = i == 10'h226 ? _GEN_2266 : _GEN_2265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2268 = io_inputBit | _GEN_2267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2269 = i == 10'h226 ? _GEN_2268 : _GEN_2267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2270 = ~io_inputBit | _GEN_2269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2271 = i == 10'h228 ? _GEN_2270 : _GEN_2269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2272 = io_inputBit ? 1'h0 : _GEN_2271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2273 = i == 10'h228 ? _GEN_2272 : _GEN_2271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2274 = ~io_inputBit ? 1'h0 : _GEN_2273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2275 = i == 10'h22a ? _GEN_2274 : _GEN_2273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2276 = io_inputBit | _GEN_2275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2277 = i == 10'h22a ? _GEN_2276 : _GEN_2275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2278 = ~io_inputBit | _GEN_2277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2279 = i == 10'h22c ? _GEN_2278 : _GEN_2277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2280 = io_inputBit ? 1'h0 : _GEN_2279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2281 = i == 10'h22c ? _GEN_2280 : _GEN_2279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2282 = ~io_inputBit ? 1'h0 : _GEN_2281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2283 = i == 10'h22e ? _GEN_2282 : _GEN_2281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2284 = io_inputBit | _GEN_2283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2285 = i == 10'h22e ? _GEN_2284 : _GEN_2283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2286 = ~io_inputBit | _GEN_2285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2287 = i == 10'h230 ? _GEN_2286 : _GEN_2285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2288 = io_inputBit ? 1'h0 : _GEN_2287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2289 = i == 10'h230 ? _GEN_2288 : _GEN_2287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2290 = ~io_inputBit ? 1'h0 : _GEN_2289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2291 = i == 10'h232 ? _GEN_2290 : _GEN_2289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2292 = io_inputBit | _GEN_2291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2293 = i == 10'h232 ? _GEN_2292 : _GEN_2291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2294 = ~io_inputBit | _GEN_2293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2295 = i == 10'h234 ? _GEN_2294 : _GEN_2293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2296 = io_inputBit ? 1'h0 : _GEN_2295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2297 = i == 10'h234 ? _GEN_2296 : _GEN_2295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2298 = ~io_inputBit ? 1'h0 : _GEN_2297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2299 = i == 10'h236 ? _GEN_2298 : _GEN_2297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2300 = io_inputBit | _GEN_2299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2301 = i == 10'h236 ? _GEN_2300 : _GEN_2299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2302 = ~io_inputBit | _GEN_2301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2303 = i == 10'h238 ? _GEN_2302 : _GEN_2301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2304 = io_inputBit ? 1'h0 : _GEN_2303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2305 = i == 10'h238 ? _GEN_2304 : _GEN_2303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2306 = ~io_inputBit ? 1'h0 : _GEN_2305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2307 = i == 10'h23a ? _GEN_2306 : _GEN_2305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2308 = io_inputBit | _GEN_2307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2309 = i == 10'h23a ? _GEN_2308 : _GEN_2307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2310 = ~io_inputBit | _GEN_2309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2311 = i == 10'h23c ? _GEN_2310 : _GEN_2309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2312 = io_inputBit ? 1'h0 : _GEN_2311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2313 = i == 10'h23c ? _GEN_2312 : _GEN_2311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2314 = ~io_inputBit ? 1'h0 : _GEN_2313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2315 = i == 10'h23e ? _GEN_2314 : _GEN_2313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2316 = io_inputBit | _GEN_2315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2317 = i == 10'h23e ? _GEN_2316 : _GEN_2315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2318 = ~io_inputBit | _GEN_2317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2319 = i == 10'h240 ? _GEN_2318 : _GEN_2317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2320 = io_inputBit ? 1'h0 : _GEN_2319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2321 = i == 10'h240 ? _GEN_2320 : _GEN_2319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2322 = ~io_inputBit ? 1'h0 : _GEN_2321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2323 = i == 10'h242 ? _GEN_2322 : _GEN_2321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2324 = io_inputBit | _GEN_2323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2325 = i == 10'h242 ? _GEN_2324 : _GEN_2323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2326 = ~io_inputBit | _GEN_2325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2327 = i == 10'h244 ? _GEN_2326 : _GEN_2325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2328 = io_inputBit ? 1'h0 : _GEN_2327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2329 = i == 10'h244 ? _GEN_2328 : _GEN_2327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2330 = ~io_inputBit ? 1'h0 : _GEN_2329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2331 = i == 10'h246 ? _GEN_2330 : _GEN_2329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2332 = io_inputBit | _GEN_2331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2333 = i == 10'h246 ? _GEN_2332 : _GEN_2331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2334 = ~io_inputBit | _GEN_2333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2335 = i == 10'h248 ? _GEN_2334 : _GEN_2333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2336 = io_inputBit ? 1'h0 : _GEN_2335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2337 = i == 10'h248 ? _GEN_2336 : _GEN_2335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2338 = io_inputBit ? 1'h0 : _GEN_1871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2339 = i == 10'h0 ? _GEN_2338 : _GEN_1871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2340 = io_inputBit ? 1'h0 : _GEN_2339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2341 = i == 10'h1 ? _GEN_2340 : _GEN_2339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2342 = io_inputBit ? 1'h0 : _GEN_2341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2343 = i == 10'h8 ? _GEN_2342 : _GEN_2341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2344 = ~io_inputBit ? 1'h0 : _GEN_2343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2345 = i == 10'hf ? _GEN_2344 : _GEN_2343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2346 = io_inputBit ? 1'h0 : _GEN_2345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2347 = i == 10'h11 ? _GEN_2346 : _GEN_2345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2348 = ~io_inputBit ? 1'h0 : _GEN_2347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2349 = i == 10'h20 ? _GEN_2348 : _GEN_2347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2350 = io_inputBit ? 1'h0 : _GEN_2349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2351 = i == 10'h48 ? _GEN_2350 : _GEN_2349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2352 = ~io_inputBit ? 1'h0 : _GEN_2351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2353 = i == 10'h10b ? _GEN_2352 : _GEN_2351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2354 = io_inputBit ? 1'h0 : _GEN_2353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2355 = i == 10'h124 ? _GEN_2354 : _GEN_2353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2356 = ~io_inputBit ? 1'h0 : _GEN_2355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2357 = i == 10'h218 ? _GEN_2356 : _GEN_2355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2358 = io_inputBit | _GEN_2357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2359 = i == 10'h218 ? _GEN_2358 : _GEN_2357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2360 = ~io_inputBit | _GEN_2359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2361 = i == 10'h219 ? _GEN_2360 : _GEN_2359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2362 = io_inputBit ? 1'h0 : _GEN_2361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2363 = i == 10'h219 ? _GEN_2362 : _GEN_2361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2364 = ~io_inputBit ? 1'h0 : _GEN_2363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2365 = i == 10'h21a ? _GEN_2364 : _GEN_2363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2366 = io_inputBit | _GEN_2365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2367 = i == 10'h21a ? _GEN_2366 : _GEN_2365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2368 = ~io_inputBit | _GEN_2367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2369 = i == 10'h21b ? _GEN_2368 : _GEN_2367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2370 = io_inputBit ? 1'h0 : _GEN_2369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2371 = i == 10'h21b ? _GEN_2370 : _GEN_2369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2372 = ~io_inputBit ? 1'h0 : _GEN_2371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2373 = i == 10'h21c ? _GEN_2372 : _GEN_2371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2374 = io_inputBit | _GEN_2373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2375 = i == 10'h21c ? _GEN_2374 : _GEN_2373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2376 = ~io_inputBit | _GEN_2375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2377 = i == 10'h21d ? _GEN_2376 : _GEN_2375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2378 = io_inputBit ? 1'h0 : _GEN_2377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2379 = i == 10'h21d ? _GEN_2378 : _GEN_2377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2380 = ~io_inputBit ? 1'h0 : _GEN_2379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2381 = i == 10'h21e ? _GEN_2380 : _GEN_2379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2382 = io_inputBit | _GEN_2381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2383 = i == 10'h21e ? _GEN_2382 : _GEN_2381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2384 = ~io_inputBit | _GEN_2383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2385 = i == 10'h21f ? _GEN_2384 : _GEN_2383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2386 = io_inputBit ? 1'h0 : _GEN_2385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2387 = i == 10'h21f ? _GEN_2386 : _GEN_2385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2388 = ~io_inputBit ? 1'h0 : _GEN_2387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2389 = i == 10'h220 ? _GEN_2388 : _GEN_2387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2390 = io_inputBit | _GEN_2389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2391 = i == 10'h220 ? _GEN_2390 : _GEN_2389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2392 = ~io_inputBit | _GEN_2391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2393 = i == 10'h221 ? _GEN_2392 : _GEN_2391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2394 = io_inputBit ? 1'h0 : _GEN_2393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2395 = i == 10'h221 ? _GEN_2394 : _GEN_2393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2396 = ~io_inputBit ? 1'h0 : _GEN_2395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2397 = i == 10'h222 ? _GEN_2396 : _GEN_2395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2398 = io_inputBit | _GEN_2397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2399 = i == 10'h222 ? _GEN_2398 : _GEN_2397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2400 = ~io_inputBit | _GEN_2399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2401 = i == 10'h223 ? _GEN_2400 : _GEN_2399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2402 = io_inputBit ? 1'h0 : _GEN_2401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2403 = i == 10'h223 ? _GEN_2402 : _GEN_2401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2404 = ~io_inputBit ? 1'h0 : _GEN_2403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2405 = i == 10'h224 ? _GEN_2404 : _GEN_2403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2406 = io_inputBit | _GEN_2405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2407 = i == 10'h224 ? _GEN_2406 : _GEN_2405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2408 = ~io_inputBit | _GEN_2407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2409 = i == 10'h225 ? _GEN_2408 : _GEN_2407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2410 = io_inputBit ? 1'h0 : _GEN_2409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2411 = i == 10'h225 ? _GEN_2410 : _GEN_2409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2412 = ~io_inputBit ? 1'h0 : _GEN_2411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2413 = i == 10'h226 ? _GEN_2412 : _GEN_2411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2414 = io_inputBit | _GEN_2413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2415 = i == 10'h226 ? _GEN_2414 : _GEN_2413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2416 = ~io_inputBit | _GEN_2415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2417 = i == 10'h227 ? _GEN_2416 : _GEN_2415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2418 = io_inputBit ? 1'h0 : _GEN_2417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2419 = i == 10'h227 ? _GEN_2418 : _GEN_2417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2420 = ~io_inputBit ? 1'h0 : _GEN_2419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2421 = i == 10'h228 ? _GEN_2420 : _GEN_2419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2422 = io_inputBit | _GEN_2421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2423 = i == 10'h228 ? _GEN_2422 : _GEN_2421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2424 = ~io_inputBit | _GEN_2423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2425 = i == 10'h229 ? _GEN_2424 : _GEN_2423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2426 = io_inputBit ? 1'h0 : _GEN_2425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2427 = i == 10'h229 ? _GEN_2426 : _GEN_2425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2428 = ~io_inputBit ? 1'h0 : _GEN_2427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2429 = i == 10'h22a ? _GEN_2428 : _GEN_2427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2430 = io_inputBit | _GEN_2429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2431 = i == 10'h22a ? _GEN_2430 : _GEN_2429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2432 = ~io_inputBit | _GEN_2431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2433 = i == 10'h22b ? _GEN_2432 : _GEN_2431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2434 = io_inputBit ? 1'h0 : _GEN_2433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2435 = i == 10'h22b ? _GEN_2434 : _GEN_2433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2436 = ~io_inputBit ? 1'h0 : _GEN_2435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2437 = i == 10'h22c ? _GEN_2436 : _GEN_2435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2438 = io_inputBit | _GEN_2437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2439 = i == 10'h22c ? _GEN_2438 : _GEN_2437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2440 = ~io_inputBit | _GEN_2439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2441 = i == 10'h22d ? _GEN_2440 : _GEN_2439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2442 = io_inputBit ? 1'h0 : _GEN_2441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2443 = i == 10'h22d ? _GEN_2442 : _GEN_2441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2444 = ~io_inputBit ? 1'h0 : _GEN_2443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2445 = i == 10'h22e ? _GEN_2444 : _GEN_2443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2446 = io_inputBit | _GEN_2445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2447 = i == 10'h22e ? _GEN_2446 : _GEN_2445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2448 = ~io_inputBit | _GEN_2447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2449 = i == 10'h22f ? _GEN_2448 : _GEN_2447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2450 = io_inputBit ? 1'h0 : _GEN_2449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2451 = i == 10'h22f ? _GEN_2450 : _GEN_2449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2452 = ~io_inputBit ? 1'h0 : _GEN_2451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2453 = i == 10'h230 ? _GEN_2452 : _GEN_2451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2454 = io_inputBit | _GEN_2453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2455 = i == 10'h230 ? _GEN_2454 : _GEN_2453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2456 = ~io_inputBit | _GEN_2455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2457 = i == 10'h231 ? _GEN_2456 : _GEN_2455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2458 = io_inputBit ? 1'h0 : _GEN_2457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2459 = i == 10'h231 ? _GEN_2458 : _GEN_2457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2460 = ~io_inputBit ? 1'h0 : _GEN_2459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2461 = i == 10'h232 ? _GEN_2460 : _GEN_2459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2462 = io_inputBit | _GEN_2461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2463 = i == 10'h232 ? _GEN_2462 : _GEN_2461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2464 = ~io_inputBit | _GEN_2463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2465 = i == 10'h233 ? _GEN_2464 : _GEN_2463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2466 = io_inputBit ? 1'h0 : _GEN_2465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2467 = i == 10'h233 ? _GEN_2466 : _GEN_2465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2468 = ~io_inputBit ? 1'h0 : _GEN_2467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2469 = i == 10'h234 ? _GEN_2468 : _GEN_2467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2470 = io_inputBit | _GEN_2469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2471 = i == 10'h234 ? _GEN_2470 : _GEN_2469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2472 = ~io_inputBit | _GEN_2471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2473 = i == 10'h235 ? _GEN_2472 : _GEN_2471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2474 = io_inputBit ? 1'h0 : _GEN_2473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2475 = i == 10'h235 ? _GEN_2474 : _GEN_2473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2476 = ~io_inputBit ? 1'h0 : _GEN_2475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2477 = i == 10'h236 ? _GEN_2476 : _GEN_2475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2478 = io_inputBit | _GEN_2477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2479 = i == 10'h236 ? _GEN_2478 : _GEN_2477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2480 = ~io_inputBit | _GEN_2479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2481 = i == 10'h237 ? _GEN_2480 : _GEN_2479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2482 = io_inputBit ? 1'h0 : _GEN_2481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2483 = i == 10'h237 ? _GEN_2482 : _GEN_2481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2484 = ~io_inputBit ? 1'h0 : _GEN_2483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2485 = i == 10'h238 ? _GEN_2484 : _GEN_2483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2486 = io_inputBit | _GEN_2485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2487 = i == 10'h238 ? _GEN_2486 : _GEN_2485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2488 = ~io_inputBit | _GEN_2487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2489 = i == 10'h239 ? _GEN_2488 : _GEN_2487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2490 = io_inputBit ? 1'h0 : _GEN_2489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2491 = i == 10'h239 ? _GEN_2490 : _GEN_2489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2492 = ~io_inputBit ? 1'h0 : _GEN_2491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2493 = i == 10'h23a ? _GEN_2492 : _GEN_2491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2494 = io_inputBit | _GEN_2493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2495 = i == 10'h23a ? _GEN_2494 : _GEN_2493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2496 = ~io_inputBit | _GEN_2495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2497 = i == 10'h23b ? _GEN_2496 : _GEN_2495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2498 = io_inputBit ? 1'h0 : _GEN_2497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2499 = i == 10'h23b ? _GEN_2498 : _GEN_2497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2500 = ~io_inputBit ? 1'h0 : _GEN_2499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2501 = i == 10'h23c ? _GEN_2500 : _GEN_2499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2502 = io_inputBit | _GEN_2501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2503 = i == 10'h23c ? _GEN_2502 : _GEN_2501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2504 = ~io_inputBit | _GEN_2503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2505 = i == 10'h23d ? _GEN_2504 : _GEN_2503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2506 = io_inputBit ? 1'h0 : _GEN_2505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2507 = i == 10'h23d ? _GEN_2506 : _GEN_2505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2508 = ~io_inputBit ? 1'h0 : _GEN_2507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2509 = i == 10'h23e ? _GEN_2508 : _GEN_2507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2510 = io_inputBit | _GEN_2509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2511 = i == 10'h23e ? _GEN_2510 : _GEN_2509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2512 = ~io_inputBit | _GEN_2511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2513 = i == 10'h23f ? _GEN_2512 : _GEN_2511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2514 = io_inputBit ? 1'h0 : _GEN_2513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2515 = i == 10'h23f ? _GEN_2514 : _GEN_2513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2516 = ~io_inputBit ? 1'h0 : _GEN_2515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2517 = i == 10'h240 ? _GEN_2516 : _GEN_2515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2518 = io_inputBit | _GEN_2517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2519 = i == 10'h240 ? _GEN_2518 : _GEN_2517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2520 = ~io_inputBit | _GEN_2519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2521 = i == 10'h241 ? _GEN_2520 : _GEN_2519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2522 = io_inputBit ? 1'h0 : _GEN_2521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2523 = i == 10'h241 ? _GEN_2522 : _GEN_2521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2524 = ~io_inputBit ? 1'h0 : _GEN_2523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2525 = i == 10'h242 ? _GEN_2524 : _GEN_2523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2526 = io_inputBit | _GEN_2525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2527 = i == 10'h242 ? _GEN_2526 : _GEN_2525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2528 = ~io_inputBit | _GEN_2527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2529 = i == 10'h243 ? _GEN_2528 : _GEN_2527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2530 = io_inputBit ? 1'h0 : _GEN_2529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2531 = i == 10'h243 ? _GEN_2530 : _GEN_2529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2532 = ~io_inputBit ? 1'h0 : _GEN_2531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2533 = i == 10'h244 ? _GEN_2532 : _GEN_2531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2534 = io_inputBit | _GEN_2533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2535 = i == 10'h244 ? _GEN_2534 : _GEN_2533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2536 = ~io_inputBit | _GEN_2535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2537 = i == 10'h245 ? _GEN_2536 : _GEN_2535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2538 = io_inputBit ? 1'h0 : _GEN_2537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2539 = i == 10'h245 ? _GEN_2538 : _GEN_2537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2540 = ~io_inputBit ? 1'h0 : _GEN_2539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2541 = i == 10'h246 ? _GEN_2540 : _GEN_2539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2542 = io_inputBit | _GEN_2541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2543 = i == 10'h246 ? _GEN_2542 : _GEN_2541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2544 = ~io_inputBit | _GEN_2543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2545 = i == 10'h247 ? _GEN_2544 : _GEN_2543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2546 = io_inputBit ? 1'h0 : _GEN_2545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2547 = i == 10'h247 ? _GEN_2546 : _GEN_2545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2548 = ~io_inputBit ? 1'h0 : _GEN_2547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2549 = i == 10'h248 ? _GEN_2548 : _GEN_2547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2550 = io_inputBit | _GEN_2549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2551 = i == 10'h248 ? _GEN_2550 : _GEN_2549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2552 = ~io_inputBit | _GEN_2551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2553 = i == 10'h249 ? _GEN_2552 : _GEN_2551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2554 = io_inputBit ? 1'h0 : _GEN_2553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2555 = i == 10'h249 ? _GEN_2554 : _GEN_2553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2556 = io_inputBit ? 1'h0 : _GEN_1921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2557 = i == 10'h0 ? _GEN_2556 : _GEN_1921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2558 = io_inputBit ? 1'h0 : _GEN_2557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2559 = i == 10'h1 ? _GEN_2558 : _GEN_2557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2560 = io_inputBit ? 1'h0 : _GEN_2559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2561 = i == 10'h8 ? _GEN_2560 : _GEN_2559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2562 = ~io_inputBit ? 1'h0 : _GEN_2561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2563 = i == 10'hf ? _GEN_2562 : _GEN_2561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2564 = io_inputBit ? 1'h0 : _GEN_2563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2565 = i == 10'h11 ? _GEN_2564 : _GEN_2563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2566 = ~io_inputBit ? 1'h0 : _GEN_2565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2567 = i == 10'h20 ? _GEN_2566 : _GEN_2565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2568 = io_inputBit ? 1'h0 : _GEN_2567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2569 = i == 10'h48 ? _GEN_2568 : _GEN_2567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2570 = ~io_inputBit ? 1'h0 : _GEN_2569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2571 = i == 10'h10b ? _GEN_2570 : _GEN_2569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2572 = io_inputBit ? 1'h0 : _GEN_2571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2573 = i == 10'h124 ? _GEN_2572 : _GEN_2571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2574 = ~io_inputBit ? 1'h0 : _GEN_2573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2575 = i == 10'h218 ? _GEN_2574 : _GEN_2573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2576 = io_inputBit | _GEN_2575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2577 = i == 10'h218 ? _GEN_2576 : _GEN_2575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2578 = ~io_inputBit ? 1'h0 : _GEN_2577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2579 = i == 10'h219 ? _GEN_2578 : _GEN_2577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2580 = io_inputBit | _GEN_2579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2581 = i == 10'h219 ? _GEN_2580 : _GEN_2579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2582 = ~io_inputBit ? 1'h0 : _GEN_2581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2583 = i == 10'h21a ? _GEN_2582 : _GEN_2581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2584 = io_inputBit | _GEN_2583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2585 = i == 10'h21a ? _GEN_2584 : _GEN_2583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2586 = ~io_inputBit ? 1'h0 : _GEN_2585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2587 = i == 10'h21b ? _GEN_2586 : _GEN_2585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2588 = io_inputBit | _GEN_2587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2589 = i == 10'h21b ? _GEN_2588 : _GEN_2587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2590 = ~io_inputBit ? 1'h0 : _GEN_2589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2591 = i == 10'h21c ? _GEN_2590 : _GEN_2589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2592 = io_inputBit | _GEN_2591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2593 = i == 10'h21c ? _GEN_2592 : _GEN_2591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2594 = ~io_inputBit ? 1'h0 : _GEN_2593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2595 = i == 10'h21d ? _GEN_2594 : _GEN_2593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2596 = io_inputBit | _GEN_2595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2597 = i == 10'h21d ? _GEN_2596 : _GEN_2595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2598 = ~io_inputBit ? 1'h0 : _GEN_2597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2599 = i == 10'h21e ? _GEN_2598 : _GEN_2597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2600 = io_inputBit | _GEN_2599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2601 = i == 10'h21e ? _GEN_2600 : _GEN_2599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2602 = ~io_inputBit ? 1'h0 : _GEN_2601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2603 = i == 10'h21f ? _GEN_2602 : _GEN_2601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2604 = io_inputBit | _GEN_2603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2605 = i == 10'h21f ? _GEN_2604 : _GEN_2603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2606 = ~io_inputBit ? 1'h0 : _GEN_2605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2607 = i == 10'h220 ? _GEN_2606 : _GEN_2605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2608 = io_inputBit | _GEN_2607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2609 = i == 10'h220 ? _GEN_2608 : _GEN_2607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2610 = ~io_inputBit ? 1'h0 : _GEN_2609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2611 = i == 10'h221 ? _GEN_2610 : _GEN_2609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2612 = io_inputBit | _GEN_2611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2613 = i == 10'h221 ? _GEN_2612 : _GEN_2611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2614 = ~io_inputBit ? 1'h0 : _GEN_2613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2615 = i == 10'h222 ? _GEN_2614 : _GEN_2613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2616 = io_inputBit | _GEN_2615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2617 = i == 10'h222 ? _GEN_2616 : _GEN_2615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2618 = ~io_inputBit ? 1'h0 : _GEN_2617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2619 = i == 10'h223 ? _GEN_2618 : _GEN_2617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2620 = io_inputBit | _GEN_2619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2621 = i == 10'h223 ? _GEN_2620 : _GEN_2619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2622 = ~io_inputBit ? 1'h0 : _GEN_2621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2623 = i == 10'h224 ? _GEN_2622 : _GEN_2621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2624 = io_inputBit | _GEN_2623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2625 = i == 10'h224 ? _GEN_2624 : _GEN_2623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2626 = ~io_inputBit ? 1'h0 : _GEN_2625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2627 = i == 10'h225 ? _GEN_2626 : _GEN_2625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2628 = io_inputBit | _GEN_2627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2629 = i == 10'h225 ? _GEN_2628 : _GEN_2627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2630 = ~io_inputBit ? 1'h0 : _GEN_2629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2631 = i == 10'h226 ? _GEN_2630 : _GEN_2629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2632 = io_inputBit | _GEN_2631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2633 = i == 10'h226 ? _GEN_2632 : _GEN_2631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2634 = ~io_inputBit ? 1'h0 : _GEN_2633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2635 = i == 10'h227 ? _GEN_2634 : _GEN_2633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2636 = io_inputBit | _GEN_2635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2637 = i == 10'h227 ? _GEN_2636 : _GEN_2635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2638 = ~io_inputBit ? 1'h0 : _GEN_2637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2639 = i == 10'h228 ? _GEN_2638 : _GEN_2637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2640 = io_inputBit | _GEN_2639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2641 = i == 10'h228 ? _GEN_2640 : _GEN_2639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2642 = ~io_inputBit ? 1'h0 : _GEN_2641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2643 = i == 10'h229 ? _GEN_2642 : _GEN_2641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2644 = io_inputBit | _GEN_2643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2645 = i == 10'h229 ? _GEN_2644 : _GEN_2643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2646 = ~io_inputBit ? 1'h0 : _GEN_2645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2647 = i == 10'h22a ? _GEN_2646 : _GEN_2645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2648 = io_inputBit | _GEN_2647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2649 = i == 10'h22a ? _GEN_2648 : _GEN_2647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2650 = ~io_inputBit ? 1'h0 : _GEN_2649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2651 = i == 10'h22b ? _GEN_2650 : _GEN_2649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2652 = io_inputBit | _GEN_2651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2653 = i == 10'h22b ? _GEN_2652 : _GEN_2651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2654 = ~io_inputBit ? 1'h0 : _GEN_2653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2655 = i == 10'h22c ? _GEN_2654 : _GEN_2653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2656 = io_inputBit | _GEN_2655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2657 = i == 10'h22c ? _GEN_2656 : _GEN_2655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2658 = ~io_inputBit ? 1'h0 : _GEN_2657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2659 = i == 10'h22d ? _GEN_2658 : _GEN_2657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2660 = io_inputBit | _GEN_2659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2661 = i == 10'h22d ? _GEN_2660 : _GEN_2659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2662 = ~io_inputBit ? 1'h0 : _GEN_2661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2663 = i == 10'h22e ? _GEN_2662 : _GEN_2661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2664 = io_inputBit | _GEN_2663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2665 = i == 10'h22e ? _GEN_2664 : _GEN_2663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2666 = ~io_inputBit ? 1'h0 : _GEN_2665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2667 = i == 10'h22f ? _GEN_2666 : _GEN_2665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2668 = io_inputBit | _GEN_2667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2669 = i == 10'h22f ? _GEN_2668 : _GEN_2667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2670 = ~io_inputBit ? 1'h0 : _GEN_2669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2671 = i == 10'h230 ? _GEN_2670 : _GEN_2669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2672 = io_inputBit | _GEN_2671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2673 = i == 10'h230 ? _GEN_2672 : _GEN_2671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2674 = ~io_inputBit ? 1'h0 : _GEN_2673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2675 = i == 10'h231 ? _GEN_2674 : _GEN_2673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2676 = io_inputBit | _GEN_2675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2677 = i == 10'h231 ? _GEN_2676 : _GEN_2675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2678 = ~io_inputBit ? 1'h0 : _GEN_2677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2679 = i == 10'h232 ? _GEN_2678 : _GEN_2677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2680 = io_inputBit | _GEN_2679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2681 = i == 10'h232 ? _GEN_2680 : _GEN_2679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2682 = ~io_inputBit ? 1'h0 : _GEN_2681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2683 = i == 10'h233 ? _GEN_2682 : _GEN_2681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2684 = io_inputBit | _GEN_2683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2685 = i == 10'h233 ? _GEN_2684 : _GEN_2683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2686 = ~io_inputBit ? 1'h0 : _GEN_2685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2687 = i == 10'h234 ? _GEN_2686 : _GEN_2685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2688 = io_inputBit | _GEN_2687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2689 = i == 10'h234 ? _GEN_2688 : _GEN_2687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2690 = ~io_inputBit ? 1'h0 : _GEN_2689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2691 = i == 10'h235 ? _GEN_2690 : _GEN_2689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2692 = io_inputBit | _GEN_2691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2693 = i == 10'h235 ? _GEN_2692 : _GEN_2691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2694 = ~io_inputBit ? 1'h0 : _GEN_2693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2695 = i == 10'h236 ? _GEN_2694 : _GEN_2693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2696 = io_inputBit | _GEN_2695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2697 = i == 10'h236 ? _GEN_2696 : _GEN_2695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2698 = ~io_inputBit ? 1'h0 : _GEN_2697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2699 = i == 10'h237 ? _GEN_2698 : _GEN_2697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2700 = io_inputBit | _GEN_2699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2701 = i == 10'h237 ? _GEN_2700 : _GEN_2699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2702 = ~io_inputBit ? 1'h0 : _GEN_2701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2703 = i == 10'h238 ? _GEN_2702 : _GEN_2701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2704 = io_inputBit | _GEN_2703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2705 = i == 10'h238 ? _GEN_2704 : _GEN_2703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2706 = ~io_inputBit ? 1'h0 : _GEN_2705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2707 = i == 10'h239 ? _GEN_2706 : _GEN_2705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2708 = io_inputBit | _GEN_2707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2709 = i == 10'h239 ? _GEN_2708 : _GEN_2707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2710 = ~io_inputBit ? 1'h0 : _GEN_2709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2711 = i == 10'h23a ? _GEN_2710 : _GEN_2709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2712 = io_inputBit | _GEN_2711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2713 = i == 10'h23a ? _GEN_2712 : _GEN_2711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2714 = ~io_inputBit ? 1'h0 : _GEN_2713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2715 = i == 10'h23b ? _GEN_2714 : _GEN_2713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2716 = io_inputBit | _GEN_2715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2717 = i == 10'h23b ? _GEN_2716 : _GEN_2715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2718 = ~io_inputBit ? 1'h0 : _GEN_2717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2719 = i == 10'h23c ? _GEN_2718 : _GEN_2717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2720 = io_inputBit | _GEN_2719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2721 = i == 10'h23c ? _GEN_2720 : _GEN_2719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2722 = ~io_inputBit ? 1'h0 : _GEN_2721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2723 = i == 10'h23d ? _GEN_2722 : _GEN_2721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2724 = io_inputBit | _GEN_2723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2725 = i == 10'h23d ? _GEN_2724 : _GEN_2723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2726 = ~io_inputBit ? 1'h0 : _GEN_2725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2727 = i == 10'h23e ? _GEN_2726 : _GEN_2725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2728 = io_inputBit | _GEN_2727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2729 = i == 10'h23e ? _GEN_2728 : _GEN_2727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2730 = ~io_inputBit ? 1'h0 : _GEN_2729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2731 = i == 10'h23f ? _GEN_2730 : _GEN_2729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2732 = io_inputBit | _GEN_2731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2733 = i == 10'h23f ? _GEN_2732 : _GEN_2731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2734 = ~io_inputBit ? 1'h0 : _GEN_2733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2735 = i == 10'h240 ? _GEN_2734 : _GEN_2733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2736 = io_inputBit | _GEN_2735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2737 = i == 10'h240 ? _GEN_2736 : _GEN_2735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2738 = ~io_inputBit ? 1'h0 : _GEN_2737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2739 = i == 10'h241 ? _GEN_2738 : _GEN_2737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2740 = io_inputBit | _GEN_2739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2741 = i == 10'h241 ? _GEN_2740 : _GEN_2739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2742 = ~io_inputBit ? 1'h0 : _GEN_2741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2743 = i == 10'h242 ? _GEN_2742 : _GEN_2741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2744 = io_inputBit | _GEN_2743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2745 = i == 10'h242 ? _GEN_2744 : _GEN_2743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2746 = ~io_inputBit ? 1'h0 : _GEN_2745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2747 = i == 10'h243 ? _GEN_2746 : _GEN_2745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2748 = io_inputBit | _GEN_2747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2749 = i == 10'h243 ? _GEN_2748 : _GEN_2747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2750 = ~io_inputBit ? 1'h0 : _GEN_2749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2751 = i == 10'h244 ? _GEN_2750 : _GEN_2749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2752 = io_inputBit | _GEN_2751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2753 = i == 10'h244 ? _GEN_2752 : _GEN_2751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2754 = ~io_inputBit ? 1'h0 : _GEN_2753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2755 = i == 10'h245 ? _GEN_2754 : _GEN_2753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2756 = io_inputBit | _GEN_2755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2757 = i == 10'h245 ? _GEN_2756 : _GEN_2755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2758 = ~io_inputBit ? 1'h0 : _GEN_2757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2759 = i == 10'h246 ? _GEN_2758 : _GEN_2757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2760 = io_inputBit | _GEN_2759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2761 = i == 10'h246 ? _GEN_2760 : _GEN_2759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2762 = ~io_inputBit ? 1'h0 : _GEN_2761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2763 = i == 10'h247 ? _GEN_2762 : _GEN_2761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2764 = io_inputBit | _GEN_2763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2765 = i == 10'h247 ? _GEN_2764 : _GEN_2763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2766 = ~io_inputBit ? 1'h0 : _GEN_2765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2767 = i == 10'h248 ? _GEN_2766 : _GEN_2765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2768 = io_inputBit | _GEN_2767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2769 = i == 10'h248 ? _GEN_2768 : _GEN_2767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2770 = ~io_inputBit ? 1'h0 : _GEN_2769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2771 = i == 10'h249 ? _GEN_2770 : _GEN_2769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2772 = io_inputBit | _GEN_2771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2773 = i == 10'h249 ? _GEN_2772 : _GEN_2771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2774 = io_inputBit ? 1'h0 : _GEN_1943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2775 = i == 10'h0 ? _GEN_2774 : _GEN_1943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2776 = io_inputBit ? 1'h0 : _GEN_2775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2777 = i == 10'h1 ? _GEN_2776 : _GEN_2775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2778 = ~io_inputBit ? 1'h0 : _GEN_2777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2779 = i == 10'h7 ? _GEN_2778 : _GEN_2777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2780 = ~io_inputBit | _GEN_2779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2781 = i == 10'h8 ? _GEN_2780 : _GEN_2779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2782 = ~io_inputBit ? 1'h0 : _GEN_2781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2783 = i == 10'h10 ? _GEN_2782 : _GEN_2781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2784 = ~io_inputBit | _GEN_2783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2785 = i == 10'h12 ? _GEN_2784 : _GEN_2783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2786 = ~io_inputBit ? 1'h0 : _GEN_2785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2787 = i == 10'h22 ? _GEN_2786 : _GEN_2785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2788 = io_inputBit ? 1'h0 : _GEN_2787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2789 = i == 10'h26 ? _GEN_2788 : _GEN_2787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2790 = io_inputBit | _GEN_2789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2791 = i == 10'h46 ? _GEN_2790 : _GEN_2789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2792 = ~io_inputBit | _GEN_2791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2793 = i == 10'h4d ? _GEN_2792 : _GEN_2791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2794 = io_inputBit | _GEN_2793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2795 = i == 10'h8d ? _GEN_2794 : _GEN_2793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2796 = ~io_inputBit | _GEN_2795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2797 = i == 10'h9c ? _GEN_2796 : _GEN_2795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2798 = ~io_inputBit ? 1'h0 : _GEN_2797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2799 = i == 10'h11b ? _GEN_2798 : _GEN_2797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2800 = io_inputBit | _GEN_2799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2801 = i == 10'h11b ? _GEN_2800 : _GEN_2799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2802 = io_inputBit ? 1'h0 : _GEN_2801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2803 = i == 10'h13a ? _GEN_2802 : _GEN_2801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2804 = ~io_inputBit | _GEN_2803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2805 = i == 10'h275 ? _GEN_2804 : _GEN_2803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2806 = io_inputBit ? 1'h0 : _GEN_2805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2807 = i == 10'h275 ? _GEN_2806 : _GEN_2805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2808 = io_inputBit ? 1'h0 : _GEN_1987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2809 = i == 10'h0 ? _GEN_2808 : _GEN_1987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2810 = io_inputBit ? 1'h0 : _GEN_2809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2811 = i == 10'h4 ? _GEN_2810 : _GEN_2809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2812 = ~io_inputBit ? 1'h0 : _GEN_2811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2813 = i == 10'h7 ? _GEN_2812 : _GEN_2811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2814 = io_inputBit ? 1'h0 : _GEN_2813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2815 = i == 10'h9 ? _GEN_2814 : _GEN_2813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2816 = io_inputBit | _GEN_2815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2817 = i == 10'h11 ? _GEN_2816 : _GEN_2815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2818 = io_inputBit ? 1'h0 : _GEN_2817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2819 = i == 10'h13 ? _GEN_2818 : _GEN_2817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2820 = ~io_inputBit ? 1'h0 : _GEN_2819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2821 = i == 10'h21 ? _GEN_2820 : _GEN_2819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2822 = ~io_inputBit | _GEN_2821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2823 = i == 10'h22 ? _GEN_2822 : _GEN_2821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2824 = ~io_inputBit ? 1'h0 : _GEN_2823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2825 = i == 10'h23 ? _GEN_2824 : _GEN_2823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2826 = io_inputBit ? 1'h0 : _GEN_2825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2827 = i == 10'h25 ? _GEN_2826 : _GEN_2825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2828 = io_inputBit | _GEN_2827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2829 = i == 10'h26 ? _GEN_2828 : _GEN_2827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2830 = io_inputBit ? 1'h0 : _GEN_2829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2831 = i == 10'h27 ? _GEN_2830 : _GEN_2829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2832 = io_inputBit | _GEN_2831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2833 = i == 10'h44 ? _GEN_2832 : _GEN_2831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2834 = io_inputBit ? 1'h0 : _GEN_2833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2835 = i == 10'h46 ? _GEN_2834 : _GEN_2833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2836 = io_inputBit | _GEN_2835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2837 = i == 10'h48 ? _GEN_2836 : _GEN_2835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2838 = ~io_inputBit | _GEN_2837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2839 = i == 10'h4b ? _GEN_2838 : _GEN_2837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2840 = ~io_inputBit ? 1'h0 : _GEN_2839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2841 = i == 10'h4d ? _GEN_2840 : _GEN_2839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2842 = ~io_inputBit | _GEN_2841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2843 = i == 10'h4f ? _GEN_2842 : _GEN_2841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2844 = io_inputBit | _GEN_2843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2845 = i == 10'h89 ? _GEN_2844 : _GEN_2843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2846 = io_inputBit ? 1'h0 : _GEN_2845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2847 = i == 10'h8d ? _GEN_2846 : _GEN_2845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2848 = io_inputBit | _GEN_2847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2849 = i == 10'h91 ? _GEN_2848 : _GEN_2847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2850 = ~io_inputBit | _GEN_2849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2851 = i == 10'h98 ? _GEN_2850 : _GEN_2849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2852 = ~io_inputBit ? 1'h0 : _GEN_2851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2853 = i == 10'h9c ? _GEN_2852 : _GEN_2851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2854 = ~io_inputBit | _GEN_2853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2855 = i == 10'ha0 ? _GEN_2854 : _GEN_2853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2856 = ~io_inputBit ? 1'h0 : _GEN_2855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2857 = i == 10'h113 ? _GEN_2856 : _GEN_2855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2858 = io_inputBit | _GEN_2857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2859 = i == 10'h113 ? _GEN_2858 : _GEN_2857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2860 = ~io_inputBit | _GEN_2859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2861 = i == 10'h11b ? _GEN_2860 : _GEN_2859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2862 = io_inputBit ? 1'h0 : _GEN_2861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2863 = i == 10'h11b ? _GEN_2862 : _GEN_2861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2864 = ~io_inputBit ? 1'h0 : _GEN_2863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2865 = i == 10'h123 ? _GEN_2864 : _GEN_2863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2866 = io_inputBit | _GEN_2865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2867 = i == 10'h123 ? _GEN_2866 : _GEN_2865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2868 = io_inputBit ? 1'h0 : _GEN_2867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2869 = i == 10'h132 ? _GEN_2868 : _GEN_2867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2870 = io_inputBit | _GEN_2869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2871 = i == 10'h13a ? _GEN_2870 : _GEN_2869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2872 = io_inputBit ? 1'h0 : _GEN_2871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2873 = i == 10'h142 ? _GEN_2872 : _GEN_2871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2874 = ~io_inputBit | _GEN_2873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2875 = i == 10'h265 ? _GEN_2874 : _GEN_2873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2876 = io_inputBit ? 1'h0 : _GEN_2875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2877 = i == 10'h265 ? _GEN_2876 : _GEN_2875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2878 = ~io_inputBit ? 1'h0 : _GEN_2877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2879 = i == 10'h275 ? _GEN_2878 : _GEN_2877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2880 = io_inputBit | _GEN_2879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2881 = i == 10'h275 ? _GEN_2880 : _GEN_2879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2882 = ~io_inputBit | _GEN_2881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2883 = i == 10'h285 ? _GEN_2882 : _GEN_2881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2884 = io_inputBit ? 1'h0 : _GEN_2883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2885 = i == 10'h285 ? _GEN_2884 : _GEN_2883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2886 = io_inputBit ? 1'h0 : _GEN_2061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2887 = i == 10'h0 ? _GEN_2886 : _GEN_2061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2888 = io_inputBit ? 1'h0 : _GEN_2887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2889 = i == 10'h4 ? _GEN_2888 : _GEN_2887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2890 = ~io_inputBit ? 1'h0 : _GEN_2889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2891 = i == 10'h7 ? _GEN_2890 : _GEN_2889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2892 = io_inputBit ? 1'h0 : _GEN_2891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2893 = i == 10'h9 ? _GEN_2892 : _GEN_2891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2894 = io_inputBit ? 1'h0 : _GEN_2893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2895 = i == 10'h11 ? _GEN_2894 : _GEN_2893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2896 = io_inputBit ? 1'h0 : _GEN_2895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2897 = i == 10'h13 ? _GEN_2896 : _GEN_2895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2898 = io_inputBit | _GEN_2897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2899 = i == 10'h43 ? _GEN_2898 : _GEN_2897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2900 = io_inputBit ? 1'h0 : _GEN_2899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2901 = i == 10'h44 ? _GEN_2900 : _GEN_2899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2902 = io_inputBit | _GEN_2901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2903 = i == 10'h45 ? _GEN_2902 : _GEN_2901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2904 = io_inputBit ? 1'h0 : _GEN_2903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2905 = i == 10'h46 ? _GEN_2904 : _GEN_2903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2906 = io_inputBit | _GEN_2905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2907 = i == 10'h47 ? _GEN_2906 : _GEN_2905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2908 = io_inputBit ? 1'h0 : _GEN_2907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2909 = i == 10'h48 ? _GEN_2908 : _GEN_2907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2910 = ~io_inputBit ? 1'h0 : _GEN_2909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2911 = i == 10'h4b ? _GEN_2910 : _GEN_2909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2912 = ~io_inputBit | _GEN_2911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2913 = i == 10'h4c ? _GEN_2912 : _GEN_2911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2914 = ~io_inputBit ? 1'h0 : _GEN_2913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2915 = i == 10'h4d ? _GEN_2914 : _GEN_2913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2916 = ~io_inputBit | _GEN_2915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2917 = i == 10'h4e ? _GEN_2916 : _GEN_2915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2918 = ~io_inputBit ? 1'h0 : _GEN_2917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2919 = i == 10'h4f ? _GEN_2918 : _GEN_2917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2920 = ~io_inputBit | _GEN_2919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2921 = i == 10'h50 ? _GEN_2920 : _GEN_2919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2922 = io_inputBit | _GEN_2921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2923 = i == 10'h87 ? _GEN_2922 : _GEN_2921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2924 = io_inputBit ? 1'h0 : _GEN_2923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2925 = i == 10'h89 ? _GEN_2924 : _GEN_2923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2926 = io_inputBit | _GEN_2925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2927 = i == 10'h8b ? _GEN_2926 : _GEN_2925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2928 = io_inputBit ? 1'h0 : _GEN_2927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2929 = i == 10'h8d ? _GEN_2928 : _GEN_2927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2930 = io_inputBit | _GEN_2929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2931 = i == 10'h8f ? _GEN_2930 : _GEN_2929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2932 = io_inputBit ? 1'h0 : _GEN_2931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2933 = i == 10'h91 ? _GEN_2932 : _GEN_2931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2934 = ~io_inputBit ? 1'h0 : _GEN_2933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2935 = i == 10'h98 ? _GEN_2934 : _GEN_2933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2936 = ~io_inputBit | _GEN_2935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2937 = i == 10'h9a ? _GEN_2936 : _GEN_2935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2938 = ~io_inputBit ? 1'h0 : _GEN_2937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2939 = i == 10'h9c ? _GEN_2938 : _GEN_2937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2940 = ~io_inputBit | _GEN_2939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2941 = i == 10'h9e ? _GEN_2940 : _GEN_2939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2942 = ~io_inputBit ? 1'h0 : _GEN_2941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2943 = i == 10'ha0 ? _GEN_2942 : _GEN_2941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2944 = ~io_inputBit | _GEN_2943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2945 = i == 10'ha2 ? _GEN_2944 : _GEN_2943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2946 = ~io_inputBit ? 1'h0 : _GEN_2945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2947 = i == 10'h10f ? _GEN_2946 : _GEN_2945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2948 = io_inputBit | _GEN_2947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2949 = i == 10'h10f ? _GEN_2948 : _GEN_2947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2950 = ~io_inputBit | _GEN_2949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2951 = i == 10'h113 ? _GEN_2950 : _GEN_2949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2952 = io_inputBit ? 1'h0 : _GEN_2951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2953 = i == 10'h113 ? _GEN_2952 : _GEN_2951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2954 = ~io_inputBit ? 1'h0 : _GEN_2953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2955 = i == 10'h117 ? _GEN_2954 : _GEN_2953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2956 = io_inputBit | _GEN_2955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2957 = i == 10'h117 ? _GEN_2956 : _GEN_2955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2958 = ~io_inputBit | _GEN_2957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2959 = i == 10'h11b ? _GEN_2958 : _GEN_2957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2960 = io_inputBit ? 1'h0 : _GEN_2959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2961 = i == 10'h11b ? _GEN_2960 : _GEN_2959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2962 = ~io_inputBit ? 1'h0 : _GEN_2961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2963 = i == 10'h11f ? _GEN_2962 : _GEN_2961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2964 = io_inputBit | _GEN_2963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2965 = i == 10'h11f ? _GEN_2964 : _GEN_2963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2966 = ~io_inputBit | _GEN_2965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2967 = i == 10'h123 ? _GEN_2966 : _GEN_2965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2968 = io_inputBit ? 1'h0 : _GEN_2967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2969 = i == 10'h123 ? _GEN_2968 : _GEN_2967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2970 = io_inputBit | _GEN_2969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2971 = i == 10'h132 ? _GEN_2970 : _GEN_2969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2972 = io_inputBit ? 1'h0 : _GEN_2971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2973 = i == 10'h136 ? _GEN_2972 : _GEN_2971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2974 = io_inputBit | _GEN_2973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2975 = i == 10'h13a ? _GEN_2974 : _GEN_2973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2976 = io_inputBit ? 1'h0 : _GEN_2975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2977 = i == 10'h13e ? _GEN_2976 : _GEN_2975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2978 = io_inputBit | _GEN_2977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2979 = i == 10'h142 ? _GEN_2978 : _GEN_2977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2980 = io_inputBit ? 1'h0 : _GEN_2979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2981 = i == 10'h146 ? _GEN_2980 : _GEN_2979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2982 = ~io_inputBit ? 1'h0 : _GEN_2981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2983 = i == 10'h265 ? _GEN_2982 : _GEN_2981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2984 = io_inputBit | _GEN_2983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2985 = i == 10'h265 ? _GEN_2984 : _GEN_2983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2986 = ~io_inputBit | _GEN_2985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2987 = i == 10'h26d ? _GEN_2986 : _GEN_2985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2988 = io_inputBit ? 1'h0 : _GEN_2987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2989 = i == 10'h26d ? _GEN_2988 : _GEN_2987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2990 = ~io_inputBit ? 1'h0 : _GEN_2989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2991 = i == 10'h275 ? _GEN_2990 : _GEN_2989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2992 = io_inputBit | _GEN_2991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2993 = i == 10'h275 ? _GEN_2992 : _GEN_2991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2994 = ~io_inputBit | _GEN_2993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2995 = i == 10'h27d ? _GEN_2994 : _GEN_2993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2996 = io_inputBit ? 1'h0 : _GEN_2995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2997 = i == 10'h27d ? _GEN_2996 : _GEN_2995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_2998 = ~io_inputBit ? 1'h0 : _GEN_2997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_2999 = i == 10'h285 ? _GEN_2998 : _GEN_2997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3000 = io_inputBit | _GEN_2999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3001 = i == 10'h285 ? _GEN_3000 : _GEN_2999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3002 = ~io_inputBit | _GEN_3001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3003 = i == 10'h28d ? _GEN_3002 : _GEN_3001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3004 = io_inputBit ? 1'h0 : _GEN_3003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3005 = i == 10'h28d ? _GEN_3004 : _GEN_3003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3006 = io_inputBit ? 1'h0 : _GEN_2171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3007 = i == 10'h0 ? _GEN_3006 : _GEN_2171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3008 = io_inputBit ? 1'h0 : _GEN_3007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3009 = i == 10'h4 ? _GEN_3008 : _GEN_3007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3010 = io_inputBit ? 1'h0 : _GEN_3009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3011 = i == 10'h9 ? _GEN_3010 : _GEN_3009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3012 = ~io_inputBit ? 1'h0 : _GEN_3011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3013 = i == 10'hf ? _GEN_3012 : _GEN_3011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3014 = io_inputBit ? 1'h0 : _GEN_3013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3015 = i == 10'h11 ? _GEN_3014 : _GEN_3013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3016 = ~io_inputBit ? 1'h0 : _GEN_3015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3017 = i == 10'h20 ? _GEN_3016 : _GEN_3015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3018 = io_inputBit ? 1'h0 : _GEN_3017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3019 = i == 10'h28 ? _GEN_3018 : _GEN_3017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3020 = ~io_inputBit ? 1'h0 : _GEN_3019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3021 = i == 10'h42 ? _GEN_3020 : _GEN_3019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3022 = io_inputBit ? 1'h0 : _GEN_3021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3023 = i == 10'h48 ? _GEN_3022 : _GEN_3021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3024 = ~io_inputBit ? 1'h0 : _GEN_3023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3025 = i == 10'h4b ? _GEN_3024 : _GEN_3023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3026 = io_inputBit ? 1'h0 : _GEN_3025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3027 = i == 10'h51 ? _GEN_3026 : _GEN_3025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3028 = io_inputBit | _GEN_3027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3029 = i == 10'h86 ? _GEN_3028 : _GEN_3027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3030 = io_inputBit ? 1'h0 : _GEN_3029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3031 = i == 10'h87 ? _GEN_3030 : _GEN_3029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3032 = io_inputBit | _GEN_3031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3033 = i == 10'h88 ? _GEN_3032 : _GEN_3031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3034 = io_inputBit ? 1'h0 : _GEN_3033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3035 = i == 10'h89 ? _GEN_3034 : _GEN_3033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3036 = io_inputBit | _GEN_3035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3037 = i == 10'h8a ? _GEN_3036 : _GEN_3035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3038 = io_inputBit ? 1'h0 : _GEN_3037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3039 = i == 10'h8b ? _GEN_3038 : _GEN_3037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3040 = io_inputBit | _GEN_3039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3041 = i == 10'h8c ? _GEN_3040 : _GEN_3039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3042 = io_inputBit ? 1'h0 : _GEN_3041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3043 = i == 10'h8d ? _GEN_3042 : _GEN_3041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3044 = io_inputBit | _GEN_3043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3045 = i == 10'h8e ? _GEN_3044 : _GEN_3043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3046 = io_inputBit ? 1'h0 : _GEN_3045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3047 = i == 10'h8f ? _GEN_3046 : _GEN_3045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3048 = io_inputBit | _GEN_3047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3049 = i == 10'h90 ? _GEN_3048 : _GEN_3047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3050 = io_inputBit ? 1'h0 : _GEN_3049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3051 = i == 10'h91 ? _GEN_3050 : _GEN_3049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3052 = ~io_inputBit ? 1'h0 : _GEN_3051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3053 = i == 10'h98 ? _GEN_3052 : _GEN_3051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3054 = ~io_inputBit | _GEN_3053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3055 = i == 10'h99 ? _GEN_3054 : _GEN_3053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3056 = ~io_inputBit ? 1'h0 : _GEN_3055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3057 = i == 10'h9a ? _GEN_3056 : _GEN_3055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3058 = ~io_inputBit | _GEN_3057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3059 = i == 10'h9b ? _GEN_3058 : _GEN_3057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3060 = ~io_inputBit ? 1'h0 : _GEN_3059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3061 = i == 10'h9c ? _GEN_3060 : _GEN_3059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3062 = ~io_inputBit | _GEN_3061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3063 = i == 10'h9d ? _GEN_3062 : _GEN_3061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3064 = ~io_inputBit ? 1'h0 : _GEN_3063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3065 = i == 10'h9e ? _GEN_3064 : _GEN_3063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3066 = ~io_inputBit | _GEN_3065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3067 = i == 10'h9f ? _GEN_3066 : _GEN_3065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3068 = ~io_inputBit ? 1'h0 : _GEN_3067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3069 = i == 10'ha0 ? _GEN_3068 : _GEN_3067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3070 = ~io_inputBit | _GEN_3069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3071 = i == 10'ha1 ? _GEN_3070 : _GEN_3069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3072 = ~io_inputBit ? 1'h0 : _GEN_3071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3073 = i == 10'ha2 ? _GEN_3072 : _GEN_3071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3074 = ~io_inputBit | _GEN_3073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3075 = i == 10'ha3 ? _GEN_3074 : _GEN_3073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3076 = ~io_inputBit ? 1'h0 : _GEN_3075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3077 = i == 10'h10d ? _GEN_3076 : _GEN_3075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3078 = io_inputBit | _GEN_3077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3079 = i == 10'h10d ? _GEN_3078 : _GEN_3077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3080 = ~io_inputBit | _GEN_3079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3081 = i == 10'h10f ? _GEN_3080 : _GEN_3079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3082 = io_inputBit ? 1'h0 : _GEN_3081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3083 = i == 10'h10f ? _GEN_3082 : _GEN_3081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3084 = ~io_inputBit ? 1'h0 : _GEN_3083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3085 = i == 10'h111 ? _GEN_3084 : _GEN_3083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3086 = io_inputBit | _GEN_3085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3087 = i == 10'h111 ? _GEN_3086 : _GEN_3085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3088 = ~io_inputBit | _GEN_3087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3089 = i == 10'h113 ? _GEN_3088 : _GEN_3087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3090 = io_inputBit ? 1'h0 : _GEN_3089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3091 = i == 10'h113 ? _GEN_3090 : _GEN_3089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3092 = ~io_inputBit ? 1'h0 : _GEN_3091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3093 = i == 10'h115 ? _GEN_3092 : _GEN_3091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3094 = io_inputBit | _GEN_3093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3095 = i == 10'h115 ? _GEN_3094 : _GEN_3093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3096 = ~io_inputBit | _GEN_3095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3097 = i == 10'h117 ? _GEN_3096 : _GEN_3095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3098 = io_inputBit ? 1'h0 : _GEN_3097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3099 = i == 10'h117 ? _GEN_3098 : _GEN_3097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3100 = ~io_inputBit ? 1'h0 : _GEN_3099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3101 = i == 10'h119 ? _GEN_3100 : _GEN_3099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3102 = io_inputBit | _GEN_3101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3103 = i == 10'h119 ? _GEN_3102 : _GEN_3101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3104 = ~io_inputBit | _GEN_3103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3105 = i == 10'h11b ? _GEN_3104 : _GEN_3103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3106 = io_inputBit ? 1'h0 : _GEN_3105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3107 = i == 10'h11b ? _GEN_3106 : _GEN_3105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3108 = ~io_inputBit ? 1'h0 : _GEN_3107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3109 = i == 10'h11d ? _GEN_3108 : _GEN_3107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3110 = io_inputBit | _GEN_3109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3111 = i == 10'h11d ? _GEN_3110 : _GEN_3109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3112 = ~io_inputBit | _GEN_3111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3113 = i == 10'h11f ? _GEN_3112 : _GEN_3111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3114 = io_inputBit ? 1'h0 : _GEN_3113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3115 = i == 10'h11f ? _GEN_3114 : _GEN_3113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3116 = ~io_inputBit ? 1'h0 : _GEN_3115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3117 = i == 10'h121 ? _GEN_3116 : _GEN_3115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3118 = io_inputBit | _GEN_3117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3119 = i == 10'h121 ? _GEN_3118 : _GEN_3117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3120 = ~io_inputBit | _GEN_3119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3121 = i == 10'h123 ? _GEN_3120 : _GEN_3119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3122 = io_inputBit ? 1'h0 : _GEN_3121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3123 = i == 10'h123 ? _GEN_3122 : _GEN_3121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3124 = io_inputBit | _GEN_3123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3125 = i == 10'h132 ? _GEN_3124 : _GEN_3123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3126 = io_inputBit ? 1'h0 : _GEN_3125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3127 = i == 10'h134 ? _GEN_3126 : _GEN_3125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3128 = io_inputBit | _GEN_3127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3129 = i == 10'h136 ? _GEN_3128 : _GEN_3127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3130 = io_inputBit ? 1'h0 : _GEN_3129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3131 = i == 10'h138 ? _GEN_3130 : _GEN_3129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3132 = io_inputBit | _GEN_3131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3133 = i == 10'h13a ? _GEN_3132 : _GEN_3131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3134 = io_inputBit ? 1'h0 : _GEN_3133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3135 = i == 10'h13c ? _GEN_3134 : _GEN_3133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3136 = io_inputBit | _GEN_3135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3137 = i == 10'h13e ? _GEN_3136 : _GEN_3135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3138 = io_inputBit ? 1'h0 : _GEN_3137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3139 = i == 10'h140 ? _GEN_3138 : _GEN_3137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3140 = io_inputBit | _GEN_3139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3141 = i == 10'h142 ? _GEN_3140 : _GEN_3139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3142 = io_inputBit ? 1'h0 : _GEN_3141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3143 = i == 10'h144 ? _GEN_3142 : _GEN_3141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3144 = io_inputBit | _GEN_3143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3145 = i == 10'h146 ? _GEN_3144 : _GEN_3143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3146 = io_inputBit ? 1'h0 : _GEN_3145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3147 = i == 10'h148 ? _GEN_3146 : _GEN_3145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3148 = ~io_inputBit ? 1'h0 : _GEN_3147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3149 = i == 10'h265 ? _GEN_3148 : _GEN_3147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3150 = io_inputBit | _GEN_3149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3151 = i == 10'h265 ? _GEN_3150 : _GEN_3149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3152 = ~io_inputBit | _GEN_3151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3153 = i == 10'h269 ? _GEN_3152 : _GEN_3151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3154 = io_inputBit ? 1'h0 : _GEN_3153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3155 = i == 10'h269 ? _GEN_3154 : _GEN_3153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3156 = ~io_inputBit ? 1'h0 : _GEN_3155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3157 = i == 10'h26d ? _GEN_3156 : _GEN_3155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3158 = io_inputBit | _GEN_3157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3159 = i == 10'h26d ? _GEN_3158 : _GEN_3157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3160 = ~io_inputBit | _GEN_3159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3161 = i == 10'h271 ? _GEN_3160 : _GEN_3159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3162 = io_inputBit ? 1'h0 : _GEN_3161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3163 = i == 10'h271 ? _GEN_3162 : _GEN_3161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3164 = ~io_inputBit ? 1'h0 : _GEN_3163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3165 = i == 10'h275 ? _GEN_3164 : _GEN_3163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3166 = io_inputBit | _GEN_3165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3167 = i == 10'h275 ? _GEN_3166 : _GEN_3165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3168 = ~io_inputBit | _GEN_3167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3169 = i == 10'h279 ? _GEN_3168 : _GEN_3167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3170 = io_inputBit ? 1'h0 : _GEN_3169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3171 = i == 10'h279 ? _GEN_3170 : _GEN_3169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3172 = ~io_inputBit ? 1'h0 : _GEN_3171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3173 = i == 10'h27d ? _GEN_3172 : _GEN_3171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3174 = io_inputBit | _GEN_3173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3175 = i == 10'h27d ? _GEN_3174 : _GEN_3173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3176 = ~io_inputBit | _GEN_3175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3177 = i == 10'h281 ? _GEN_3176 : _GEN_3175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3178 = io_inputBit ? 1'h0 : _GEN_3177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3179 = i == 10'h281 ? _GEN_3178 : _GEN_3177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3180 = ~io_inputBit ? 1'h0 : _GEN_3179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3181 = i == 10'h285 ? _GEN_3180 : _GEN_3179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3182 = io_inputBit | _GEN_3181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3183 = i == 10'h285 ? _GEN_3182 : _GEN_3181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3184 = ~io_inputBit | _GEN_3183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3185 = i == 10'h289 ? _GEN_3184 : _GEN_3183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3186 = io_inputBit ? 1'h0 : _GEN_3185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3187 = i == 10'h289 ? _GEN_3186 : _GEN_3185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3188 = ~io_inputBit ? 1'h0 : _GEN_3187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3189 = i == 10'h28d ? _GEN_3188 : _GEN_3187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3190 = io_inputBit | _GEN_3189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3191 = i == 10'h28d ? _GEN_3190 : _GEN_3189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3192 = ~io_inputBit | _GEN_3191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3193 = i == 10'h291 ? _GEN_3192 : _GEN_3191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3194 = io_inputBit ? 1'h0 : _GEN_3193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3195 = i == 10'h291 ? _GEN_3194 : _GEN_3193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3196 = io_inputBit ? 1'h0 : _GEN_2337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3197 = i == 10'h0 ? _GEN_3196 : _GEN_2337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3198 = io_inputBit ? 1'h0 : _GEN_3197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3199 = i == 10'h4 ? _GEN_3198 : _GEN_3197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3200 = io_inputBit ? 1'h0 : _GEN_3199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3201 = i == 10'h9 ? _GEN_3200 : _GEN_3199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3202 = ~io_inputBit ? 1'h0 : _GEN_3201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3203 = i == 10'hf ? _GEN_3202 : _GEN_3201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3204 = io_inputBit | _GEN_3203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3205 = i == 10'h11 ? _GEN_3204 : _GEN_3203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3206 = ~io_inputBit ? 1'h0 : _GEN_3205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3207 = i == 10'h20 ? _GEN_3206 : _GEN_3205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3208 = io_inputBit ? 1'h0 : _GEN_3207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3209 = i == 10'h28 ? _GEN_3208 : _GEN_3207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3210 = io_inputBit | _GEN_3209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3211 = i == 10'h48 ? _GEN_3210 : _GEN_3209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3212 = ~io_inputBit | _GEN_3211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3213 = i == 10'h4b ? _GEN_3212 : _GEN_3211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3214 = ~io_inputBit ? 1'h0 : _GEN_3213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3215 = i == 10'h85 ? _GEN_3214 : _GEN_3213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3216 = io_inputBit ? 1'h0 : _GEN_3215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3217 = i == 10'ha4 ? _GEN_3216 : _GEN_3215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3218 = ~io_inputBit ? 1'h0 : _GEN_3217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3219 = i == 10'h10c ? _GEN_3218 : _GEN_3217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3220 = io_inputBit | _GEN_3219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3221 = i == 10'h10c ? _GEN_3220 : _GEN_3219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3222 = ~io_inputBit | _GEN_3221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3223 = i == 10'h10d ? _GEN_3222 : _GEN_3221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3224 = io_inputBit ? 1'h0 : _GEN_3223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3225 = i == 10'h10d ? _GEN_3224 : _GEN_3223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3226 = ~io_inputBit ? 1'h0 : _GEN_3225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3227 = i == 10'h10e ? _GEN_3226 : _GEN_3225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3228 = io_inputBit | _GEN_3227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3229 = i == 10'h10e ? _GEN_3228 : _GEN_3227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3230 = ~io_inputBit | _GEN_3229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3231 = i == 10'h10f ? _GEN_3230 : _GEN_3229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3232 = io_inputBit ? 1'h0 : _GEN_3231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3233 = i == 10'h10f ? _GEN_3232 : _GEN_3231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3234 = ~io_inputBit ? 1'h0 : _GEN_3233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3235 = i == 10'h110 ? _GEN_3234 : _GEN_3233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3236 = io_inputBit | _GEN_3235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3237 = i == 10'h110 ? _GEN_3236 : _GEN_3235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3238 = ~io_inputBit | _GEN_3237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3239 = i == 10'h111 ? _GEN_3238 : _GEN_3237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3240 = io_inputBit ? 1'h0 : _GEN_3239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3241 = i == 10'h111 ? _GEN_3240 : _GEN_3239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3242 = ~io_inputBit ? 1'h0 : _GEN_3241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3243 = i == 10'h112 ? _GEN_3242 : _GEN_3241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3244 = io_inputBit | _GEN_3243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3245 = i == 10'h112 ? _GEN_3244 : _GEN_3243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3246 = ~io_inputBit | _GEN_3245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3247 = i == 10'h113 ? _GEN_3246 : _GEN_3245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3248 = io_inputBit ? 1'h0 : _GEN_3247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3249 = i == 10'h113 ? _GEN_3248 : _GEN_3247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3250 = ~io_inputBit ? 1'h0 : _GEN_3249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3251 = i == 10'h114 ? _GEN_3250 : _GEN_3249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3252 = io_inputBit | _GEN_3251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3253 = i == 10'h114 ? _GEN_3252 : _GEN_3251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3254 = ~io_inputBit | _GEN_3253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3255 = i == 10'h115 ? _GEN_3254 : _GEN_3253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3256 = io_inputBit ? 1'h0 : _GEN_3255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3257 = i == 10'h115 ? _GEN_3256 : _GEN_3255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3258 = ~io_inputBit ? 1'h0 : _GEN_3257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3259 = i == 10'h116 ? _GEN_3258 : _GEN_3257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3260 = io_inputBit | _GEN_3259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3261 = i == 10'h116 ? _GEN_3260 : _GEN_3259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3262 = ~io_inputBit | _GEN_3261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3263 = i == 10'h117 ? _GEN_3262 : _GEN_3261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3264 = io_inputBit ? 1'h0 : _GEN_3263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3265 = i == 10'h117 ? _GEN_3264 : _GEN_3263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3266 = ~io_inputBit ? 1'h0 : _GEN_3265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3267 = i == 10'h118 ? _GEN_3266 : _GEN_3265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3268 = io_inputBit | _GEN_3267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3269 = i == 10'h118 ? _GEN_3268 : _GEN_3267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3270 = ~io_inputBit | _GEN_3269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3271 = i == 10'h119 ? _GEN_3270 : _GEN_3269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3272 = io_inputBit ? 1'h0 : _GEN_3271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3273 = i == 10'h119 ? _GEN_3272 : _GEN_3271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3274 = ~io_inputBit ? 1'h0 : _GEN_3273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3275 = i == 10'h11a ? _GEN_3274 : _GEN_3273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3276 = io_inputBit | _GEN_3275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3277 = i == 10'h11a ? _GEN_3276 : _GEN_3275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3278 = ~io_inputBit | _GEN_3277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3279 = i == 10'h11b ? _GEN_3278 : _GEN_3277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3280 = io_inputBit ? 1'h0 : _GEN_3279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3281 = i == 10'h11b ? _GEN_3280 : _GEN_3279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3282 = ~io_inputBit ? 1'h0 : _GEN_3281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3283 = i == 10'h11c ? _GEN_3282 : _GEN_3281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3284 = io_inputBit | _GEN_3283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3285 = i == 10'h11c ? _GEN_3284 : _GEN_3283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3286 = ~io_inputBit | _GEN_3285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3287 = i == 10'h11d ? _GEN_3286 : _GEN_3285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3288 = io_inputBit ? 1'h0 : _GEN_3287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3289 = i == 10'h11d ? _GEN_3288 : _GEN_3287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3290 = ~io_inputBit ? 1'h0 : _GEN_3289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3291 = i == 10'h11e ? _GEN_3290 : _GEN_3289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3292 = io_inputBit | _GEN_3291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3293 = i == 10'h11e ? _GEN_3292 : _GEN_3291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3294 = ~io_inputBit | _GEN_3293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3295 = i == 10'h11f ? _GEN_3294 : _GEN_3293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3296 = io_inputBit ? 1'h0 : _GEN_3295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3297 = i == 10'h11f ? _GEN_3296 : _GEN_3295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3298 = ~io_inputBit ? 1'h0 : _GEN_3297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3299 = i == 10'h120 ? _GEN_3298 : _GEN_3297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3300 = io_inputBit | _GEN_3299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3301 = i == 10'h120 ? _GEN_3300 : _GEN_3299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3302 = ~io_inputBit | _GEN_3301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3303 = i == 10'h121 ? _GEN_3302 : _GEN_3301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3304 = io_inputBit ? 1'h0 : _GEN_3303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3305 = i == 10'h121 ? _GEN_3304 : _GEN_3303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3306 = ~io_inputBit ? 1'h0 : _GEN_3305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3307 = i == 10'h122 ? _GEN_3306 : _GEN_3305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3308 = io_inputBit | _GEN_3307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3309 = i == 10'h122 ? _GEN_3308 : _GEN_3307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3310 = ~io_inputBit | _GEN_3309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3311 = i == 10'h123 ? _GEN_3310 : _GEN_3309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3312 = io_inputBit ? 1'h0 : _GEN_3311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3313 = i == 10'h123 ? _GEN_3312 : _GEN_3311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3314 = ~io_inputBit ? 1'h0 : _GEN_3313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3315 = i == 10'h124 ? _GEN_3314 : _GEN_3313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3316 = io_inputBit | _GEN_3315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3317 = i == 10'h124 ? _GEN_3316 : _GEN_3315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3318 = io_inputBit ? 1'h0 : _GEN_3317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3319 = i == 10'h131 ? _GEN_3318 : _GEN_3317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3320 = io_inputBit | _GEN_3319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3321 = i == 10'h132 ? _GEN_3320 : _GEN_3319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3322 = io_inputBit ? 1'h0 : _GEN_3321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3323 = i == 10'h133 ? _GEN_3322 : _GEN_3321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3324 = io_inputBit | _GEN_3323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3325 = i == 10'h134 ? _GEN_3324 : _GEN_3323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3326 = io_inputBit ? 1'h0 : _GEN_3325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3327 = i == 10'h135 ? _GEN_3326 : _GEN_3325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3328 = io_inputBit | _GEN_3327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3329 = i == 10'h136 ? _GEN_3328 : _GEN_3327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3330 = io_inputBit ? 1'h0 : _GEN_3329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3331 = i == 10'h137 ? _GEN_3330 : _GEN_3329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3332 = io_inputBit | _GEN_3331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3333 = i == 10'h138 ? _GEN_3332 : _GEN_3331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3334 = io_inputBit ? 1'h0 : _GEN_3333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3335 = i == 10'h139 ? _GEN_3334 : _GEN_3333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3336 = io_inputBit | _GEN_3335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3337 = i == 10'h13a ? _GEN_3336 : _GEN_3335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3338 = io_inputBit ? 1'h0 : _GEN_3337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3339 = i == 10'h13b ? _GEN_3338 : _GEN_3337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3340 = io_inputBit | _GEN_3339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3341 = i == 10'h13c ? _GEN_3340 : _GEN_3339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3342 = io_inputBit ? 1'h0 : _GEN_3341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3343 = i == 10'h13d ? _GEN_3342 : _GEN_3341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3344 = io_inputBit | _GEN_3343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3345 = i == 10'h13e ? _GEN_3344 : _GEN_3343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3346 = io_inputBit ? 1'h0 : _GEN_3345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3347 = i == 10'h13f ? _GEN_3346 : _GEN_3345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3348 = io_inputBit | _GEN_3347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3349 = i == 10'h140 ? _GEN_3348 : _GEN_3347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3350 = io_inputBit ? 1'h0 : _GEN_3349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3351 = i == 10'h141 ? _GEN_3350 : _GEN_3349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3352 = io_inputBit | _GEN_3351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3353 = i == 10'h142 ? _GEN_3352 : _GEN_3351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3354 = io_inputBit ? 1'h0 : _GEN_3353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3355 = i == 10'h143 ? _GEN_3354 : _GEN_3353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3356 = io_inputBit | _GEN_3355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3357 = i == 10'h144 ? _GEN_3356 : _GEN_3355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3358 = io_inputBit ? 1'h0 : _GEN_3357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3359 = i == 10'h145 ? _GEN_3358 : _GEN_3357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3360 = io_inputBit | _GEN_3359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3361 = i == 10'h146 ? _GEN_3360 : _GEN_3359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3362 = io_inputBit ? 1'h0 : _GEN_3361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3363 = i == 10'h147 ? _GEN_3362 : _GEN_3361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3364 = io_inputBit | _GEN_3363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3365 = i == 10'h148 ? _GEN_3364 : _GEN_3363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3366 = io_inputBit ? 1'h0 : _GEN_3365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3367 = i == 10'h149 ? _GEN_3366 : _GEN_3365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3368 = ~io_inputBit | _GEN_3367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3369 = i == 10'h263 ? _GEN_3368 : _GEN_3367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3370 = io_inputBit ? 1'h0 : _GEN_3369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3371 = i == 10'h263 ? _GEN_3370 : _GEN_3369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3372 = ~io_inputBit ? 1'h0 : _GEN_3371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3373 = i == 10'h265 ? _GEN_3372 : _GEN_3371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3374 = io_inputBit | _GEN_3373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3375 = i == 10'h265 ? _GEN_3374 : _GEN_3373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3376 = ~io_inputBit | _GEN_3375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3377 = i == 10'h267 ? _GEN_3376 : _GEN_3375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3378 = io_inputBit ? 1'h0 : _GEN_3377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3379 = i == 10'h267 ? _GEN_3378 : _GEN_3377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3380 = ~io_inputBit ? 1'h0 : _GEN_3379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3381 = i == 10'h269 ? _GEN_3380 : _GEN_3379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3382 = io_inputBit | _GEN_3381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3383 = i == 10'h269 ? _GEN_3382 : _GEN_3381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3384 = ~io_inputBit | _GEN_3383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3385 = i == 10'h26b ? _GEN_3384 : _GEN_3383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3386 = io_inputBit ? 1'h0 : _GEN_3385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3387 = i == 10'h26b ? _GEN_3386 : _GEN_3385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3388 = ~io_inputBit ? 1'h0 : _GEN_3387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3389 = i == 10'h26d ? _GEN_3388 : _GEN_3387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3390 = io_inputBit | _GEN_3389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3391 = i == 10'h26d ? _GEN_3390 : _GEN_3389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3392 = ~io_inputBit | _GEN_3391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3393 = i == 10'h26f ? _GEN_3392 : _GEN_3391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3394 = io_inputBit ? 1'h0 : _GEN_3393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3395 = i == 10'h26f ? _GEN_3394 : _GEN_3393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3396 = ~io_inputBit ? 1'h0 : _GEN_3395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3397 = i == 10'h271 ? _GEN_3396 : _GEN_3395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3398 = io_inputBit | _GEN_3397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3399 = i == 10'h271 ? _GEN_3398 : _GEN_3397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3400 = ~io_inputBit | _GEN_3399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3401 = i == 10'h273 ? _GEN_3400 : _GEN_3399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3402 = io_inputBit ? 1'h0 : _GEN_3401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3403 = i == 10'h273 ? _GEN_3402 : _GEN_3401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3404 = ~io_inputBit ? 1'h0 : _GEN_3403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3405 = i == 10'h275 ? _GEN_3404 : _GEN_3403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3406 = io_inputBit | _GEN_3405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3407 = i == 10'h275 ? _GEN_3406 : _GEN_3405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3408 = ~io_inputBit | _GEN_3407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3409 = i == 10'h277 ? _GEN_3408 : _GEN_3407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3410 = io_inputBit ? 1'h0 : _GEN_3409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3411 = i == 10'h277 ? _GEN_3410 : _GEN_3409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3412 = ~io_inputBit ? 1'h0 : _GEN_3411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3413 = i == 10'h279 ? _GEN_3412 : _GEN_3411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3414 = io_inputBit | _GEN_3413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3415 = i == 10'h279 ? _GEN_3414 : _GEN_3413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3416 = ~io_inputBit | _GEN_3415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3417 = i == 10'h27b ? _GEN_3416 : _GEN_3415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3418 = io_inputBit ? 1'h0 : _GEN_3417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3419 = i == 10'h27b ? _GEN_3418 : _GEN_3417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3420 = ~io_inputBit ? 1'h0 : _GEN_3419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3421 = i == 10'h27d ? _GEN_3420 : _GEN_3419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3422 = io_inputBit | _GEN_3421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3423 = i == 10'h27d ? _GEN_3422 : _GEN_3421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3424 = ~io_inputBit | _GEN_3423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3425 = i == 10'h27f ? _GEN_3424 : _GEN_3423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3426 = io_inputBit ? 1'h0 : _GEN_3425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3427 = i == 10'h27f ? _GEN_3426 : _GEN_3425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3428 = ~io_inputBit ? 1'h0 : _GEN_3427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3429 = i == 10'h281 ? _GEN_3428 : _GEN_3427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3430 = io_inputBit | _GEN_3429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3431 = i == 10'h281 ? _GEN_3430 : _GEN_3429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3432 = ~io_inputBit | _GEN_3431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3433 = i == 10'h283 ? _GEN_3432 : _GEN_3431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3434 = io_inputBit ? 1'h0 : _GEN_3433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3435 = i == 10'h283 ? _GEN_3434 : _GEN_3433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3436 = ~io_inputBit ? 1'h0 : _GEN_3435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3437 = i == 10'h285 ? _GEN_3436 : _GEN_3435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3438 = io_inputBit | _GEN_3437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3439 = i == 10'h285 ? _GEN_3438 : _GEN_3437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3440 = ~io_inputBit | _GEN_3439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3441 = i == 10'h287 ? _GEN_3440 : _GEN_3439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3442 = io_inputBit ? 1'h0 : _GEN_3441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3443 = i == 10'h287 ? _GEN_3442 : _GEN_3441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3444 = ~io_inputBit ? 1'h0 : _GEN_3443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3445 = i == 10'h289 ? _GEN_3444 : _GEN_3443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3446 = io_inputBit | _GEN_3445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3447 = i == 10'h289 ? _GEN_3446 : _GEN_3445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3448 = ~io_inputBit | _GEN_3447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3449 = i == 10'h28b ? _GEN_3448 : _GEN_3447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3450 = io_inputBit ? 1'h0 : _GEN_3449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3451 = i == 10'h28b ? _GEN_3450 : _GEN_3449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3452 = ~io_inputBit ? 1'h0 : _GEN_3451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3453 = i == 10'h28d ? _GEN_3452 : _GEN_3451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3454 = io_inputBit | _GEN_3453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3455 = i == 10'h28d ? _GEN_3454 : _GEN_3453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3456 = ~io_inputBit | _GEN_3455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3457 = i == 10'h28f ? _GEN_3456 : _GEN_3455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3458 = io_inputBit ? 1'h0 : _GEN_3457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3459 = i == 10'h28f ? _GEN_3458 : _GEN_3457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3460 = ~io_inputBit ? 1'h0 : _GEN_3459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3461 = i == 10'h291 ? _GEN_3460 : _GEN_3459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3462 = io_inputBit | _GEN_3461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3463 = i == 10'h291 ? _GEN_3462 : _GEN_3461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3464 = ~io_inputBit | _GEN_3463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3465 = i == 10'h293 ? _GEN_3464 : _GEN_3463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3466 = io_inputBit ? 1'h0 : _GEN_3465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3467 = i == 10'h293 ? _GEN_3466 : _GEN_3465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3468 = io_inputBit ? 1'h0 : _GEN_2555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3469 = i == 10'h0 ? _GEN_3468 : _GEN_2555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3470 = io_inputBit ? 1'h0 : _GEN_3469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3471 = i == 10'h4 ? _GEN_3470 : _GEN_3469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3472 = io_inputBit ? 1'h0 : _GEN_3471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3473 = i == 10'h9 ? _GEN_3472 : _GEN_3471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3474 = ~io_inputBit ? 1'h0 : _GEN_3473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3475 = i == 10'hf ? _GEN_3474 : _GEN_3473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3476 = io_inputBit ? 1'h0 : _GEN_3475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3477 = i == 10'h11 ? _GEN_3476 : _GEN_3475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3478 = ~io_inputBit ? 1'h0 : _GEN_3477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3479 = i == 10'h20 ? _GEN_3478 : _GEN_3477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3480 = io_inputBit ? 1'h0 : _GEN_3479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3481 = i == 10'h28 ? _GEN_3480 : _GEN_3479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3482 = io_inputBit ? 1'h0 : _GEN_3481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3483 = i == 10'h48 ? _GEN_3482 : _GEN_3481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3484 = ~io_inputBit ? 1'h0 : _GEN_3483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3485 = i == 10'h4b ? _GEN_3484 : _GEN_3483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3486 = ~io_inputBit ? 1'h0 : _GEN_3485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3487 = i == 10'h85 ? _GEN_3486 : _GEN_3485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3488 = io_inputBit ? 1'h0 : _GEN_3487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3489 = i == 10'ha4 ? _GEN_3488 : _GEN_3487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3490 = ~io_inputBit | _GEN_3489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3491 = i == 10'h10c ? _GEN_3490 : _GEN_3489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3492 = io_inputBit ? 1'h0 : _GEN_3491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3493 = i == 10'h10c ? _GEN_3492 : _GEN_3491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3494 = ~io_inputBit | _GEN_3493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3495 = i == 10'h10d ? _GEN_3494 : _GEN_3493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3496 = io_inputBit ? 1'h0 : _GEN_3495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3497 = i == 10'h10d ? _GEN_3496 : _GEN_3495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3498 = ~io_inputBit | _GEN_3497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3499 = i == 10'h10e ? _GEN_3498 : _GEN_3497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3500 = io_inputBit ? 1'h0 : _GEN_3499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3501 = i == 10'h10e ? _GEN_3500 : _GEN_3499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3502 = ~io_inputBit | _GEN_3501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3503 = i == 10'h10f ? _GEN_3502 : _GEN_3501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3504 = io_inputBit ? 1'h0 : _GEN_3503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3505 = i == 10'h10f ? _GEN_3504 : _GEN_3503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3506 = ~io_inputBit | _GEN_3505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3507 = i == 10'h110 ? _GEN_3506 : _GEN_3505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3508 = io_inputBit ? 1'h0 : _GEN_3507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3509 = i == 10'h110 ? _GEN_3508 : _GEN_3507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3510 = ~io_inputBit | _GEN_3509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3511 = i == 10'h111 ? _GEN_3510 : _GEN_3509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3512 = io_inputBit ? 1'h0 : _GEN_3511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3513 = i == 10'h111 ? _GEN_3512 : _GEN_3511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3514 = ~io_inputBit | _GEN_3513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3515 = i == 10'h112 ? _GEN_3514 : _GEN_3513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3516 = io_inputBit ? 1'h0 : _GEN_3515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3517 = i == 10'h112 ? _GEN_3516 : _GEN_3515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3518 = ~io_inputBit | _GEN_3517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3519 = i == 10'h113 ? _GEN_3518 : _GEN_3517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3520 = io_inputBit ? 1'h0 : _GEN_3519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3521 = i == 10'h113 ? _GEN_3520 : _GEN_3519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3522 = ~io_inputBit | _GEN_3521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3523 = i == 10'h114 ? _GEN_3522 : _GEN_3521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3524 = io_inputBit ? 1'h0 : _GEN_3523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3525 = i == 10'h114 ? _GEN_3524 : _GEN_3523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3526 = ~io_inputBit | _GEN_3525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3527 = i == 10'h115 ? _GEN_3526 : _GEN_3525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3528 = io_inputBit ? 1'h0 : _GEN_3527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3529 = i == 10'h115 ? _GEN_3528 : _GEN_3527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3530 = ~io_inputBit | _GEN_3529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3531 = i == 10'h116 ? _GEN_3530 : _GEN_3529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3532 = io_inputBit ? 1'h0 : _GEN_3531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3533 = i == 10'h116 ? _GEN_3532 : _GEN_3531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3534 = ~io_inputBit | _GEN_3533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3535 = i == 10'h117 ? _GEN_3534 : _GEN_3533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3536 = io_inputBit ? 1'h0 : _GEN_3535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3537 = i == 10'h117 ? _GEN_3536 : _GEN_3535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3538 = ~io_inputBit | _GEN_3537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3539 = i == 10'h118 ? _GEN_3538 : _GEN_3537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3540 = io_inputBit ? 1'h0 : _GEN_3539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3541 = i == 10'h118 ? _GEN_3540 : _GEN_3539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3542 = ~io_inputBit | _GEN_3541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3543 = i == 10'h119 ? _GEN_3542 : _GEN_3541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3544 = io_inputBit ? 1'h0 : _GEN_3543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3545 = i == 10'h119 ? _GEN_3544 : _GEN_3543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3546 = ~io_inputBit | _GEN_3545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3547 = i == 10'h11a ? _GEN_3546 : _GEN_3545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3548 = io_inputBit ? 1'h0 : _GEN_3547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3549 = i == 10'h11a ? _GEN_3548 : _GEN_3547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3550 = ~io_inputBit | _GEN_3549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3551 = i == 10'h11b ? _GEN_3550 : _GEN_3549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3552 = io_inputBit ? 1'h0 : _GEN_3551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3553 = i == 10'h11b ? _GEN_3552 : _GEN_3551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3554 = ~io_inputBit | _GEN_3553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3555 = i == 10'h11c ? _GEN_3554 : _GEN_3553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3556 = io_inputBit ? 1'h0 : _GEN_3555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3557 = i == 10'h11c ? _GEN_3556 : _GEN_3555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3558 = ~io_inputBit | _GEN_3557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3559 = i == 10'h11d ? _GEN_3558 : _GEN_3557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3560 = io_inputBit ? 1'h0 : _GEN_3559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3561 = i == 10'h11d ? _GEN_3560 : _GEN_3559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3562 = ~io_inputBit | _GEN_3561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3563 = i == 10'h11e ? _GEN_3562 : _GEN_3561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3564 = io_inputBit ? 1'h0 : _GEN_3563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3565 = i == 10'h11e ? _GEN_3564 : _GEN_3563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3566 = ~io_inputBit | _GEN_3565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3567 = i == 10'h11f ? _GEN_3566 : _GEN_3565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3568 = io_inputBit ? 1'h0 : _GEN_3567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3569 = i == 10'h11f ? _GEN_3568 : _GEN_3567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3570 = ~io_inputBit | _GEN_3569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3571 = i == 10'h120 ? _GEN_3570 : _GEN_3569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3572 = io_inputBit ? 1'h0 : _GEN_3571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3573 = i == 10'h120 ? _GEN_3572 : _GEN_3571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3574 = ~io_inputBit | _GEN_3573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3575 = i == 10'h121 ? _GEN_3574 : _GEN_3573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3576 = io_inputBit ? 1'h0 : _GEN_3575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3577 = i == 10'h121 ? _GEN_3576 : _GEN_3575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3578 = ~io_inputBit | _GEN_3577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3579 = i == 10'h122 ? _GEN_3578 : _GEN_3577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3580 = io_inputBit ? 1'h0 : _GEN_3579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3581 = i == 10'h122 ? _GEN_3580 : _GEN_3579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3582 = ~io_inputBit | _GEN_3581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3583 = i == 10'h123 ? _GEN_3582 : _GEN_3581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3584 = io_inputBit ? 1'h0 : _GEN_3583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3585 = i == 10'h123 ? _GEN_3584 : _GEN_3583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3586 = ~io_inputBit | _GEN_3585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3587 = i == 10'h124 ? _GEN_3586 : _GEN_3585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3588 = io_inputBit ? 1'h0 : _GEN_3587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3589 = i == 10'h124 ? _GEN_3588 : _GEN_3587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3590 = ~io_inputBit ? 1'h0 : _GEN_3589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3591 = i == 10'h263 ? _GEN_3590 : _GEN_3589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3592 = io_inputBit | _GEN_3591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3593 = i == 10'h263 ? _GEN_3592 : _GEN_3591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3594 = ~io_inputBit | _GEN_3593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3595 = i == 10'h264 ? _GEN_3594 : _GEN_3593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3596 = io_inputBit ? 1'h0 : _GEN_3595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3597 = i == 10'h264 ? _GEN_3596 : _GEN_3595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3598 = ~io_inputBit ? 1'h0 : _GEN_3597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3599 = i == 10'h265 ? _GEN_3598 : _GEN_3597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3600 = io_inputBit | _GEN_3599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3601 = i == 10'h265 ? _GEN_3600 : _GEN_3599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3602 = ~io_inputBit | _GEN_3601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3603 = i == 10'h266 ? _GEN_3602 : _GEN_3601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3604 = io_inputBit ? 1'h0 : _GEN_3603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3605 = i == 10'h266 ? _GEN_3604 : _GEN_3603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3606 = ~io_inputBit ? 1'h0 : _GEN_3605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3607 = i == 10'h267 ? _GEN_3606 : _GEN_3605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3608 = io_inputBit | _GEN_3607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3609 = i == 10'h267 ? _GEN_3608 : _GEN_3607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3610 = ~io_inputBit | _GEN_3609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3611 = i == 10'h268 ? _GEN_3610 : _GEN_3609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3612 = io_inputBit ? 1'h0 : _GEN_3611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3613 = i == 10'h268 ? _GEN_3612 : _GEN_3611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3614 = ~io_inputBit ? 1'h0 : _GEN_3613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3615 = i == 10'h269 ? _GEN_3614 : _GEN_3613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3616 = io_inputBit | _GEN_3615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3617 = i == 10'h269 ? _GEN_3616 : _GEN_3615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3618 = ~io_inputBit | _GEN_3617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3619 = i == 10'h26a ? _GEN_3618 : _GEN_3617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3620 = io_inputBit ? 1'h0 : _GEN_3619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3621 = i == 10'h26a ? _GEN_3620 : _GEN_3619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3622 = ~io_inputBit ? 1'h0 : _GEN_3621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3623 = i == 10'h26b ? _GEN_3622 : _GEN_3621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3624 = io_inputBit | _GEN_3623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3625 = i == 10'h26b ? _GEN_3624 : _GEN_3623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3626 = ~io_inputBit | _GEN_3625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3627 = i == 10'h26c ? _GEN_3626 : _GEN_3625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3628 = io_inputBit ? 1'h0 : _GEN_3627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3629 = i == 10'h26c ? _GEN_3628 : _GEN_3627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3630 = ~io_inputBit ? 1'h0 : _GEN_3629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3631 = i == 10'h26d ? _GEN_3630 : _GEN_3629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3632 = io_inputBit | _GEN_3631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3633 = i == 10'h26d ? _GEN_3632 : _GEN_3631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3634 = ~io_inputBit | _GEN_3633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3635 = i == 10'h26e ? _GEN_3634 : _GEN_3633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3636 = io_inputBit ? 1'h0 : _GEN_3635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3637 = i == 10'h26e ? _GEN_3636 : _GEN_3635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3638 = ~io_inputBit ? 1'h0 : _GEN_3637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3639 = i == 10'h26f ? _GEN_3638 : _GEN_3637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3640 = io_inputBit | _GEN_3639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3641 = i == 10'h26f ? _GEN_3640 : _GEN_3639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3642 = ~io_inputBit | _GEN_3641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3643 = i == 10'h270 ? _GEN_3642 : _GEN_3641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3644 = io_inputBit ? 1'h0 : _GEN_3643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3645 = i == 10'h270 ? _GEN_3644 : _GEN_3643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3646 = ~io_inputBit ? 1'h0 : _GEN_3645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3647 = i == 10'h271 ? _GEN_3646 : _GEN_3645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3648 = io_inputBit | _GEN_3647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3649 = i == 10'h271 ? _GEN_3648 : _GEN_3647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3650 = ~io_inputBit | _GEN_3649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3651 = i == 10'h272 ? _GEN_3650 : _GEN_3649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3652 = io_inputBit ? 1'h0 : _GEN_3651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3653 = i == 10'h272 ? _GEN_3652 : _GEN_3651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3654 = ~io_inputBit ? 1'h0 : _GEN_3653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3655 = i == 10'h273 ? _GEN_3654 : _GEN_3653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3656 = io_inputBit | _GEN_3655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3657 = i == 10'h273 ? _GEN_3656 : _GEN_3655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3658 = ~io_inputBit | _GEN_3657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3659 = i == 10'h274 ? _GEN_3658 : _GEN_3657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3660 = io_inputBit ? 1'h0 : _GEN_3659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3661 = i == 10'h274 ? _GEN_3660 : _GEN_3659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3662 = ~io_inputBit ? 1'h0 : _GEN_3661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3663 = i == 10'h275 ? _GEN_3662 : _GEN_3661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3664 = io_inputBit | _GEN_3663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3665 = i == 10'h275 ? _GEN_3664 : _GEN_3663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3666 = ~io_inputBit | _GEN_3665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3667 = i == 10'h276 ? _GEN_3666 : _GEN_3665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3668 = io_inputBit ? 1'h0 : _GEN_3667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3669 = i == 10'h276 ? _GEN_3668 : _GEN_3667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3670 = ~io_inputBit ? 1'h0 : _GEN_3669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3671 = i == 10'h277 ? _GEN_3670 : _GEN_3669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3672 = io_inputBit | _GEN_3671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3673 = i == 10'h277 ? _GEN_3672 : _GEN_3671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3674 = ~io_inputBit | _GEN_3673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3675 = i == 10'h278 ? _GEN_3674 : _GEN_3673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3676 = io_inputBit ? 1'h0 : _GEN_3675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3677 = i == 10'h278 ? _GEN_3676 : _GEN_3675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3678 = ~io_inputBit ? 1'h0 : _GEN_3677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3679 = i == 10'h279 ? _GEN_3678 : _GEN_3677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3680 = io_inputBit | _GEN_3679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3681 = i == 10'h279 ? _GEN_3680 : _GEN_3679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3682 = ~io_inputBit | _GEN_3681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3683 = i == 10'h27a ? _GEN_3682 : _GEN_3681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3684 = io_inputBit ? 1'h0 : _GEN_3683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3685 = i == 10'h27a ? _GEN_3684 : _GEN_3683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3686 = ~io_inputBit ? 1'h0 : _GEN_3685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3687 = i == 10'h27b ? _GEN_3686 : _GEN_3685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3688 = io_inputBit | _GEN_3687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3689 = i == 10'h27b ? _GEN_3688 : _GEN_3687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3690 = ~io_inputBit | _GEN_3689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3691 = i == 10'h27c ? _GEN_3690 : _GEN_3689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3692 = io_inputBit ? 1'h0 : _GEN_3691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3693 = i == 10'h27c ? _GEN_3692 : _GEN_3691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3694 = ~io_inputBit ? 1'h0 : _GEN_3693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3695 = i == 10'h27d ? _GEN_3694 : _GEN_3693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3696 = io_inputBit | _GEN_3695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3697 = i == 10'h27d ? _GEN_3696 : _GEN_3695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3698 = ~io_inputBit | _GEN_3697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3699 = i == 10'h27e ? _GEN_3698 : _GEN_3697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3700 = io_inputBit ? 1'h0 : _GEN_3699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3701 = i == 10'h27e ? _GEN_3700 : _GEN_3699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3702 = ~io_inputBit ? 1'h0 : _GEN_3701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3703 = i == 10'h27f ? _GEN_3702 : _GEN_3701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3704 = io_inputBit | _GEN_3703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3705 = i == 10'h27f ? _GEN_3704 : _GEN_3703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3706 = ~io_inputBit | _GEN_3705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3707 = i == 10'h280 ? _GEN_3706 : _GEN_3705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3708 = io_inputBit ? 1'h0 : _GEN_3707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3709 = i == 10'h280 ? _GEN_3708 : _GEN_3707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3710 = ~io_inputBit ? 1'h0 : _GEN_3709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3711 = i == 10'h281 ? _GEN_3710 : _GEN_3709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3712 = io_inputBit | _GEN_3711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3713 = i == 10'h281 ? _GEN_3712 : _GEN_3711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3714 = ~io_inputBit | _GEN_3713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3715 = i == 10'h282 ? _GEN_3714 : _GEN_3713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3716 = io_inputBit ? 1'h0 : _GEN_3715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3717 = i == 10'h282 ? _GEN_3716 : _GEN_3715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3718 = ~io_inputBit ? 1'h0 : _GEN_3717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3719 = i == 10'h283 ? _GEN_3718 : _GEN_3717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3720 = io_inputBit | _GEN_3719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3721 = i == 10'h283 ? _GEN_3720 : _GEN_3719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3722 = ~io_inputBit | _GEN_3721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3723 = i == 10'h284 ? _GEN_3722 : _GEN_3721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3724 = io_inputBit ? 1'h0 : _GEN_3723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3725 = i == 10'h284 ? _GEN_3724 : _GEN_3723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3726 = ~io_inputBit ? 1'h0 : _GEN_3725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3727 = i == 10'h285 ? _GEN_3726 : _GEN_3725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3728 = io_inputBit | _GEN_3727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3729 = i == 10'h285 ? _GEN_3728 : _GEN_3727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3730 = ~io_inputBit | _GEN_3729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3731 = i == 10'h286 ? _GEN_3730 : _GEN_3729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3732 = io_inputBit ? 1'h0 : _GEN_3731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3733 = i == 10'h286 ? _GEN_3732 : _GEN_3731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3734 = ~io_inputBit ? 1'h0 : _GEN_3733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3735 = i == 10'h287 ? _GEN_3734 : _GEN_3733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3736 = io_inputBit | _GEN_3735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3737 = i == 10'h287 ? _GEN_3736 : _GEN_3735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3738 = ~io_inputBit | _GEN_3737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3739 = i == 10'h288 ? _GEN_3738 : _GEN_3737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3740 = io_inputBit ? 1'h0 : _GEN_3739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3741 = i == 10'h288 ? _GEN_3740 : _GEN_3739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3742 = ~io_inputBit ? 1'h0 : _GEN_3741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3743 = i == 10'h289 ? _GEN_3742 : _GEN_3741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3744 = io_inputBit | _GEN_3743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3745 = i == 10'h289 ? _GEN_3744 : _GEN_3743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3746 = ~io_inputBit | _GEN_3745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3747 = i == 10'h28a ? _GEN_3746 : _GEN_3745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3748 = io_inputBit ? 1'h0 : _GEN_3747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3749 = i == 10'h28a ? _GEN_3748 : _GEN_3747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3750 = ~io_inputBit ? 1'h0 : _GEN_3749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3751 = i == 10'h28b ? _GEN_3750 : _GEN_3749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3752 = io_inputBit | _GEN_3751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3753 = i == 10'h28b ? _GEN_3752 : _GEN_3751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3754 = ~io_inputBit | _GEN_3753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3755 = i == 10'h28c ? _GEN_3754 : _GEN_3753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3756 = io_inputBit ? 1'h0 : _GEN_3755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3757 = i == 10'h28c ? _GEN_3756 : _GEN_3755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3758 = ~io_inputBit ? 1'h0 : _GEN_3757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3759 = i == 10'h28d ? _GEN_3758 : _GEN_3757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3760 = io_inputBit | _GEN_3759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3761 = i == 10'h28d ? _GEN_3760 : _GEN_3759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3762 = ~io_inputBit | _GEN_3761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3763 = i == 10'h28e ? _GEN_3762 : _GEN_3761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3764 = io_inputBit ? 1'h0 : _GEN_3763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3765 = i == 10'h28e ? _GEN_3764 : _GEN_3763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3766 = ~io_inputBit ? 1'h0 : _GEN_3765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3767 = i == 10'h28f ? _GEN_3766 : _GEN_3765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3768 = io_inputBit | _GEN_3767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3769 = i == 10'h28f ? _GEN_3768 : _GEN_3767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3770 = ~io_inputBit | _GEN_3769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3771 = i == 10'h290 ? _GEN_3770 : _GEN_3769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3772 = io_inputBit ? 1'h0 : _GEN_3771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3773 = i == 10'h290 ? _GEN_3772 : _GEN_3771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3774 = ~io_inputBit ? 1'h0 : _GEN_3773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3775 = i == 10'h291 ? _GEN_3774 : _GEN_3773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3776 = io_inputBit | _GEN_3775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3777 = i == 10'h291 ? _GEN_3776 : _GEN_3775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3778 = ~io_inputBit | _GEN_3777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3779 = i == 10'h292 ? _GEN_3778 : _GEN_3777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3780 = io_inputBit ? 1'h0 : _GEN_3779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3781 = i == 10'h292 ? _GEN_3780 : _GEN_3779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3782 = ~io_inputBit ? 1'h0 : _GEN_3781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3783 = i == 10'h293 ? _GEN_3782 : _GEN_3781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3784 = io_inputBit | _GEN_3783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3785 = i == 10'h293 ? _GEN_3784 : _GEN_3783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3786 = ~io_inputBit | _GEN_3785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3787 = i == 10'h294 ? _GEN_3786 : _GEN_3785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3788 = io_inputBit ? 1'h0 : _GEN_3787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3789 = i == 10'h294 ? _GEN_3788 : _GEN_3787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3790 = io_inputBit ? 1'h0 : _GEN_2773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3791 = i == 10'h0 ? _GEN_3790 : _GEN_2773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3792 = io_inputBit ? 1'h0 : _GEN_3791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3793 = i == 10'h4 ? _GEN_3792 : _GEN_3791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3794 = io_inputBit ? 1'h0 : _GEN_3793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3795 = i == 10'h9 ? _GEN_3794 : _GEN_3793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3796 = ~io_inputBit ? 1'h0 : _GEN_3795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3797 = i == 10'hf ? _GEN_3796 : _GEN_3795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3798 = io_inputBit ? 1'h0 : _GEN_3797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3799 = i == 10'h11 ? _GEN_3798 : _GEN_3797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3800 = ~io_inputBit ? 1'h0 : _GEN_3799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3801 = i == 10'h20 ? _GEN_3800 : _GEN_3799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3802 = io_inputBit ? 1'h0 : _GEN_3801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3803 = i == 10'h28 ? _GEN_3802 : _GEN_3801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3804 = io_inputBit ? 1'h0 : _GEN_3803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3805 = i == 10'h48 ? _GEN_3804 : _GEN_3803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3806 = ~io_inputBit ? 1'h0 : _GEN_3805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3807 = i == 10'h4b ? _GEN_3806 : _GEN_3805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3808 = io_inputBit ? 1'h0 : _GEN_3807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3809 = i == 10'ha4 ? _GEN_3808 : _GEN_3807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3810 = ~io_inputBit ? 1'h0 : _GEN_3809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3811 = i == 10'h10b ? _GEN_3810 : _GEN_3809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3812 = io_inputBit ? 1'h0 : _GEN_3811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3813 = i == 10'h124 ? _GEN_3812 : _GEN_3811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3814 = ~io_inputBit ? 1'h0 : _GEN_3813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3815 = i == 10'h218 ? _GEN_3814 : _GEN_3813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3816 = io_inputBit | _GEN_3815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3817 = i == 10'h218 ? _GEN_3816 : _GEN_3815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3818 = ~io_inputBit ? 1'h0 : _GEN_3817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3819 = i == 10'h219 ? _GEN_3818 : _GEN_3817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3820 = io_inputBit | _GEN_3819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3821 = i == 10'h219 ? _GEN_3820 : _GEN_3819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3822 = ~io_inputBit ? 1'h0 : _GEN_3821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3823 = i == 10'h21a ? _GEN_3822 : _GEN_3821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3824 = io_inputBit | _GEN_3823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3825 = i == 10'h21a ? _GEN_3824 : _GEN_3823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3826 = ~io_inputBit ? 1'h0 : _GEN_3825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3827 = i == 10'h21b ? _GEN_3826 : _GEN_3825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3828 = io_inputBit | _GEN_3827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3829 = i == 10'h21b ? _GEN_3828 : _GEN_3827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3830 = ~io_inputBit ? 1'h0 : _GEN_3829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3831 = i == 10'h21c ? _GEN_3830 : _GEN_3829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3832 = io_inputBit | _GEN_3831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3833 = i == 10'h21c ? _GEN_3832 : _GEN_3831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3834 = ~io_inputBit ? 1'h0 : _GEN_3833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3835 = i == 10'h21d ? _GEN_3834 : _GEN_3833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3836 = io_inputBit | _GEN_3835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3837 = i == 10'h21d ? _GEN_3836 : _GEN_3835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3838 = ~io_inputBit ? 1'h0 : _GEN_3837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3839 = i == 10'h21e ? _GEN_3838 : _GEN_3837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3840 = io_inputBit | _GEN_3839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3841 = i == 10'h21e ? _GEN_3840 : _GEN_3839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3842 = ~io_inputBit ? 1'h0 : _GEN_3841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3843 = i == 10'h21f ? _GEN_3842 : _GEN_3841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3844 = io_inputBit | _GEN_3843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3845 = i == 10'h21f ? _GEN_3844 : _GEN_3843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3846 = ~io_inputBit ? 1'h0 : _GEN_3845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3847 = i == 10'h220 ? _GEN_3846 : _GEN_3845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3848 = io_inputBit | _GEN_3847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3849 = i == 10'h220 ? _GEN_3848 : _GEN_3847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3850 = ~io_inputBit ? 1'h0 : _GEN_3849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3851 = i == 10'h221 ? _GEN_3850 : _GEN_3849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3852 = io_inputBit | _GEN_3851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3853 = i == 10'h221 ? _GEN_3852 : _GEN_3851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3854 = ~io_inputBit ? 1'h0 : _GEN_3853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3855 = i == 10'h222 ? _GEN_3854 : _GEN_3853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3856 = io_inputBit | _GEN_3855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3857 = i == 10'h222 ? _GEN_3856 : _GEN_3855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3858 = ~io_inputBit ? 1'h0 : _GEN_3857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3859 = i == 10'h223 ? _GEN_3858 : _GEN_3857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3860 = io_inputBit | _GEN_3859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3861 = i == 10'h223 ? _GEN_3860 : _GEN_3859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3862 = ~io_inputBit ? 1'h0 : _GEN_3861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3863 = i == 10'h224 ? _GEN_3862 : _GEN_3861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3864 = io_inputBit | _GEN_3863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3865 = i == 10'h224 ? _GEN_3864 : _GEN_3863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3866 = ~io_inputBit ? 1'h0 : _GEN_3865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3867 = i == 10'h225 ? _GEN_3866 : _GEN_3865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3868 = io_inputBit | _GEN_3867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3869 = i == 10'h225 ? _GEN_3868 : _GEN_3867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3870 = ~io_inputBit ? 1'h0 : _GEN_3869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3871 = i == 10'h226 ? _GEN_3870 : _GEN_3869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3872 = io_inputBit | _GEN_3871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3873 = i == 10'h226 ? _GEN_3872 : _GEN_3871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3874 = ~io_inputBit ? 1'h0 : _GEN_3873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3875 = i == 10'h227 ? _GEN_3874 : _GEN_3873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3876 = io_inputBit | _GEN_3875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3877 = i == 10'h227 ? _GEN_3876 : _GEN_3875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3878 = ~io_inputBit ? 1'h0 : _GEN_3877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3879 = i == 10'h228 ? _GEN_3878 : _GEN_3877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3880 = io_inputBit | _GEN_3879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3881 = i == 10'h228 ? _GEN_3880 : _GEN_3879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3882 = ~io_inputBit ? 1'h0 : _GEN_3881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3883 = i == 10'h229 ? _GEN_3882 : _GEN_3881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3884 = io_inputBit | _GEN_3883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3885 = i == 10'h229 ? _GEN_3884 : _GEN_3883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3886 = ~io_inputBit ? 1'h0 : _GEN_3885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3887 = i == 10'h22a ? _GEN_3886 : _GEN_3885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3888 = io_inputBit | _GEN_3887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3889 = i == 10'h22a ? _GEN_3888 : _GEN_3887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3890 = ~io_inputBit ? 1'h0 : _GEN_3889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3891 = i == 10'h22b ? _GEN_3890 : _GEN_3889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3892 = io_inputBit | _GEN_3891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3893 = i == 10'h22b ? _GEN_3892 : _GEN_3891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3894 = ~io_inputBit ? 1'h0 : _GEN_3893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3895 = i == 10'h22c ? _GEN_3894 : _GEN_3893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3896 = io_inputBit | _GEN_3895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3897 = i == 10'h22c ? _GEN_3896 : _GEN_3895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3898 = ~io_inputBit ? 1'h0 : _GEN_3897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3899 = i == 10'h22d ? _GEN_3898 : _GEN_3897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3900 = io_inputBit | _GEN_3899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3901 = i == 10'h22d ? _GEN_3900 : _GEN_3899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3902 = ~io_inputBit ? 1'h0 : _GEN_3901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3903 = i == 10'h22e ? _GEN_3902 : _GEN_3901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3904 = io_inputBit | _GEN_3903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3905 = i == 10'h22e ? _GEN_3904 : _GEN_3903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3906 = ~io_inputBit ? 1'h0 : _GEN_3905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3907 = i == 10'h22f ? _GEN_3906 : _GEN_3905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3908 = io_inputBit | _GEN_3907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3909 = i == 10'h22f ? _GEN_3908 : _GEN_3907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3910 = ~io_inputBit ? 1'h0 : _GEN_3909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3911 = i == 10'h230 ? _GEN_3910 : _GEN_3909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3912 = io_inputBit | _GEN_3911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3913 = i == 10'h230 ? _GEN_3912 : _GEN_3911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3914 = ~io_inputBit ? 1'h0 : _GEN_3913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3915 = i == 10'h231 ? _GEN_3914 : _GEN_3913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3916 = io_inputBit | _GEN_3915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3917 = i == 10'h231 ? _GEN_3916 : _GEN_3915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3918 = ~io_inputBit ? 1'h0 : _GEN_3917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3919 = i == 10'h232 ? _GEN_3918 : _GEN_3917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3920 = io_inputBit | _GEN_3919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3921 = i == 10'h232 ? _GEN_3920 : _GEN_3919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3922 = ~io_inputBit ? 1'h0 : _GEN_3921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3923 = i == 10'h233 ? _GEN_3922 : _GEN_3921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3924 = io_inputBit | _GEN_3923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3925 = i == 10'h233 ? _GEN_3924 : _GEN_3923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3926 = ~io_inputBit ? 1'h0 : _GEN_3925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3927 = i == 10'h234 ? _GEN_3926 : _GEN_3925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3928 = io_inputBit | _GEN_3927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3929 = i == 10'h234 ? _GEN_3928 : _GEN_3927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3930 = ~io_inputBit ? 1'h0 : _GEN_3929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3931 = i == 10'h235 ? _GEN_3930 : _GEN_3929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3932 = io_inputBit | _GEN_3931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3933 = i == 10'h235 ? _GEN_3932 : _GEN_3931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3934 = ~io_inputBit ? 1'h0 : _GEN_3933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3935 = i == 10'h236 ? _GEN_3934 : _GEN_3933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3936 = io_inputBit | _GEN_3935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3937 = i == 10'h236 ? _GEN_3936 : _GEN_3935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3938 = ~io_inputBit ? 1'h0 : _GEN_3937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3939 = i == 10'h237 ? _GEN_3938 : _GEN_3937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3940 = io_inputBit | _GEN_3939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3941 = i == 10'h237 ? _GEN_3940 : _GEN_3939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3942 = ~io_inputBit ? 1'h0 : _GEN_3941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3943 = i == 10'h238 ? _GEN_3942 : _GEN_3941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3944 = io_inputBit | _GEN_3943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3945 = i == 10'h238 ? _GEN_3944 : _GEN_3943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3946 = ~io_inputBit ? 1'h0 : _GEN_3945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3947 = i == 10'h239 ? _GEN_3946 : _GEN_3945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3948 = io_inputBit | _GEN_3947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3949 = i == 10'h239 ? _GEN_3948 : _GEN_3947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3950 = ~io_inputBit ? 1'h0 : _GEN_3949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3951 = i == 10'h23a ? _GEN_3950 : _GEN_3949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3952 = io_inputBit | _GEN_3951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3953 = i == 10'h23a ? _GEN_3952 : _GEN_3951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3954 = ~io_inputBit ? 1'h0 : _GEN_3953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3955 = i == 10'h23b ? _GEN_3954 : _GEN_3953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3956 = io_inputBit | _GEN_3955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3957 = i == 10'h23b ? _GEN_3956 : _GEN_3955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3958 = ~io_inputBit ? 1'h0 : _GEN_3957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3959 = i == 10'h23c ? _GEN_3958 : _GEN_3957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3960 = io_inputBit | _GEN_3959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3961 = i == 10'h23c ? _GEN_3960 : _GEN_3959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3962 = ~io_inputBit ? 1'h0 : _GEN_3961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3963 = i == 10'h23d ? _GEN_3962 : _GEN_3961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3964 = io_inputBit | _GEN_3963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3965 = i == 10'h23d ? _GEN_3964 : _GEN_3963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3966 = ~io_inputBit ? 1'h0 : _GEN_3965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3967 = i == 10'h23e ? _GEN_3966 : _GEN_3965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3968 = io_inputBit | _GEN_3967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3969 = i == 10'h23e ? _GEN_3968 : _GEN_3967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3970 = ~io_inputBit ? 1'h0 : _GEN_3969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3971 = i == 10'h23f ? _GEN_3970 : _GEN_3969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3972 = io_inputBit | _GEN_3971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3973 = i == 10'h23f ? _GEN_3972 : _GEN_3971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3974 = ~io_inputBit ? 1'h0 : _GEN_3973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3975 = i == 10'h240 ? _GEN_3974 : _GEN_3973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3976 = io_inputBit | _GEN_3975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3977 = i == 10'h240 ? _GEN_3976 : _GEN_3975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3978 = ~io_inputBit ? 1'h0 : _GEN_3977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3979 = i == 10'h241 ? _GEN_3978 : _GEN_3977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3980 = io_inputBit | _GEN_3979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3981 = i == 10'h241 ? _GEN_3980 : _GEN_3979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3982 = ~io_inputBit ? 1'h0 : _GEN_3981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3983 = i == 10'h242 ? _GEN_3982 : _GEN_3981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3984 = io_inputBit | _GEN_3983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3985 = i == 10'h242 ? _GEN_3984 : _GEN_3983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3986 = ~io_inputBit ? 1'h0 : _GEN_3985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3987 = i == 10'h243 ? _GEN_3986 : _GEN_3985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3988 = io_inputBit | _GEN_3987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3989 = i == 10'h243 ? _GEN_3988 : _GEN_3987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3990 = ~io_inputBit ? 1'h0 : _GEN_3989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3991 = i == 10'h244 ? _GEN_3990 : _GEN_3989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3992 = io_inputBit | _GEN_3991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3993 = i == 10'h244 ? _GEN_3992 : _GEN_3991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3994 = ~io_inputBit ? 1'h0 : _GEN_3993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3995 = i == 10'h245 ? _GEN_3994 : _GEN_3993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3996 = io_inputBit | _GEN_3995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3997 = i == 10'h245 ? _GEN_3996 : _GEN_3995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_3998 = ~io_inputBit ? 1'h0 : _GEN_3997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3999 = i == 10'h246 ? _GEN_3998 : _GEN_3997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4000 = io_inputBit | _GEN_3999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4001 = i == 10'h246 ? _GEN_4000 : _GEN_3999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4002 = ~io_inputBit ? 1'h0 : _GEN_4001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4003 = i == 10'h247 ? _GEN_4002 : _GEN_4001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4004 = io_inputBit | _GEN_4003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4005 = i == 10'h247 ? _GEN_4004 : _GEN_4003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4006 = ~io_inputBit ? 1'h0 : _GEN_4005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4007 = i == 10'h248 ? _GEN_4006 : _GEN_4005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4008 = io_inputBit | _GEN_4007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4009 = i == 10'h248 ? _GEN_4008 : _GEN_4007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4010 = ~io_inputBit ? 1'h0 : _GEN_4009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4011 = i == 10'h249 ? _GEN_4010 : _GEN_4009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4012 = io_inputBit | _GEN_4011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4013 = i == 10'h249 ? _GEN_4012 : _GEN_4011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4014 = ~io_inputBit ? 1'h0 : _GEN_4013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4015 = i == 10'h263 ? _GEN_4014 : _GEN_4013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4016 = io_inputBit | _GEN_4015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4017 = i == 10'h263 ? _GEN_4016 : _GEN_4015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4018 = ~io_inputBit ? 1'h0 : _GEN_4017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4019 = i == 10'h264 ? _GEN_4018 : _GEN_4017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4020 = io_inputBit | _GEN_4019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4021 = i == 10'h264 ? _GEN_4020 : _GEN_4019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4022 = ~io_inputBit ? 1'h0 : _GEN_4021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4023 = i == 10'h265 ? _GEN_4022 : _GEN_4021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4024 = io_inputBit | _GEN_4023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4025 = i == 10'h265 ? _GEN_4024 : _GEN_4023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4026 = ~io_inputBit ? 1'h0 : _GEN_4025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4027 = i == 10'h266 ? _GEN_4026 : _GEN_4025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4028 = io_inputBit | _GEN_4027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4029 = i == 10'h266 ? _GEN_4028 : _GEN_4027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4030 = ~io_inputBit ? 1'h0 : _GEN_4029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4031 = i == 10'h267 ? _GEN_4030 : _GEN_4029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4032 = io_inputBit | _GEN_4031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4033 = i == 10'h267 ? _GEN_4032 : _GEN_4031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4034 = ~io_inputBit ? 1'h0 : _GEN_4033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4035 = i == 10'h268 ? _GEN_4034 : _GEN_4033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4036 = io_inputBit | _GEN_4035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4037 = i == 10'h268 ? _GEN_4036 : _GEN_4035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4038 = ~io_inputBit ? 1'h0 : _GEN_4037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4039 = i == 10'h269 ? _GEN_4038 : _GEN_4037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4040 = io_inputBit | _GEN_4039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4041 = i == 10'h269 ? _GEN_4040 : _GEN_4039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4042 = ~io_inputBit ? 1'h0 : _GEN_4041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4043 = i == 10'h26a ? _GEN_4042 : _GEN_4041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4044 = io_inputBit | _GEN_4043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4045 = i == 10'h26a ? _GEN_4044 : _GEN_4043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4046 = ~io_inputBit ? 1'h0 : _GEN_4045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4047 = i == 10'h26b ? _GEN_4046 : _GEN_4045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4048 = io_inputBit | _GEN_4047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4049 = i == 10'h26b ? _GEN_4048 : _GEN_4047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4050 = ~io_inputBit ? 1'h0 : _GEN_4049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4051 = i == 10'h26c ? _GEN_4050 : _GEN_4049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4052 = io_inputBit | _GEN_4051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4053 = i == 10'h26c ? _GEN_4052 : _GEN_4051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4054 = ~io_inputBit ? 1'h0 : _GEN_4053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4055 = i == 10'h26d ? _GEN_4054 : _GEN_4053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4056 = io_inputBit | _GEN_4055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4057 = i == 10'h26d ? _GEN_4056 : _GEN_4055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4058 = ~io_inputBit ? 1'h0 : _GEN_4057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4059 = i == 10'h26e ? _GEN_4058 : _GEN_4057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4060 = io_inputBit | _GEN_4059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4061 = i == 10'h26e ? _GEN_4060 : _GEN_4059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4062 = ~io_inputBit ? 1'h0 : _GEN_4061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4063 = i == 10'h26f ? _GEN_4062 : _GEN_4061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4064 = io_inputBit | _GEN_4063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4065 = i == 10'h26f ? _GEN_4064 : _GEN_4063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4066 = ~io_inputBit ? 1'h0 : _GEN_4065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4067 = i == 10'h270 ? _GEN_4066 : _GEN_4065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4068 = io_inputBit | _GEN_4067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4069 = i == 10'h270 ? _GEN_4068 : _GEN_4067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4070 = ~io_inputBit ? 1'h0 : _GEN_4069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4071 = i == 10'h271 ? _GEN_4070 : _GEN_4069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4072 = io_inputBit | _GEN_4071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4073 = i == 10'h271 ? _GEN_4072 : _GEN_4071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4074 = ~io_inputBit ? 1'h0 : _GEN_4073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4075 = i == 10'h272 ? _GEN_4074 : _GEN_4073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4076 = io_inputBit | _GEN_4075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4077 = i == 10'h272 ? _GEN_4076 : _GEN_4075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4078 = ~io_inputBit ? 1'h0 : _GEN_4077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4079 = i == 10'h273 ? _GEN_4078 : _GEN_4077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4080 = io_inputBit | _GEN_4079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4081 = i == 10'h273 ? _GEN_4080 : _GEN_4079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4082 = ~io_inputBit ? 1'h0 : _GEN_4081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4083 = i == 10'h274 ? _GEN_4082 : _GEN_4081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4084 = io_inputBit | _GEN_4083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4085 = i == 10'h274 ? _GEN_4084 : _GEN_4083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4086 = ~io_inputBit ? 1'h0 : _GEN_4085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4087 = i == 10'h275 ? _GEN_4086 : _GEN_4085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4088 = io_inputBit | _GEN_4087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4089 = i == 10'h275 ? _GEN_4088 : _GEN_4087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4090 = ~io_inputBit ? 1'h0 : _GEN_4089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4091 = i == 10'h276 ? _GEN_4090 : _GEN_4089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4092 = io_inputBit | _GEN_4091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4093 = i == 10'h276 ? _GEN_4092 : _GEN_4091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4094 = ~io_inputBit ? 1'h0 : _GEN_4093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4095 = i == 10'h277 ? _GEN_4094 : _GEN_4093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4096 = io_inputBit | _GEN_4095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4097 = i == 10'h277 ? _GEN_4096 : _GEN_4095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4098 = ~io_inputBit ? 1'h0 : _GEN_4097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4099 = i == 10'h278 ? _GEN_4098 : _GEN_4097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4100 = io_inputBit | _GEN_4099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4101 = i == 10'h278 ? _GEN_4100 : _GEN_4099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4102 = ~io_inputBit ? 1'h0 : _GEN_4101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4103 = i == 10'h279 ? _GEN_4102 : _GEN_4101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4104 = io_inputBit | _GEN_4103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4105 = i == 10'h279 ? _GEN_4104 : _GEN_4103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4106 = ~io_inputBit ? 1'h0 : _GEN_4105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4107 = i == 10'h27a ? _GEN_4106 : _GEN_4105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4108 = io_inputBit | _GEN_4107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4109 = i == 10'h27a ? _GEN_4108 : _GEN_4107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4110 = ~io_inputBit ? 1'h0 : _GEN_4109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4111 = i == 10'h27b ? _GEN_4110 : _GEN_4109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4112 = io_inputBit | _GEN_4111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4113 = i == 10'h27b ? _GEN_4112 : _GEN_4111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4114 = ~io_inputBit ? 1'h0 : _GEN_4113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4115 = i == 10'h27c ? _GEN_4114 : _GEN_4113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4116 = io_inputBit | _GEN_4115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4117 = i == 10'h27c ? _GEN_4116 : _GEN_4115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4118 = ~io_inputBit ? 1'h0 : _GEN_4117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4119 = i == 10'h27d ? _GEN_4118 : _GEN_4117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4120 = io_inputBit | _GEN_4119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4121 = i == 10'h27d ? _GEN_4120 : _GEN_4119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4122 = ~io_inputBit ? 1'h0 : _GEN_4121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4123 = i == 10'h27e ? _GEN_4122 : _GEN_4121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4124 = io_inputBit | _GEN_4123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4125 = i == 10'h27e ? _GEN_4124 : _GEN_4123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4126 = ~io_inputBit ? 1'h0 : _GEN_4125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4127 = i == 10'h27f ? _GEN_4126 : _GEN_4125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4128 = io_inputBit | _GEN_4127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4129 = i == 10'h27f ? _GEN_4128 : _GEN_4127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4130 = ~io_inputBit ? 1'h0 : _GEN_4129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4131 = i == 10'h280 ? _GEN_4130 : _GEN_4129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4132 = io_inputBit | _GEN_4131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4133 = i == 10'h280 ? _GEN_4132 : _GEN_4131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4134 = ~io_inputBit ? 1'h0 : _GEN_4133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4135 = i == 10'h281 ? _GEN_4134 : _GEN_4133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4136 = io_inputBit | _GEN_4135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4137 = i == 10'h281 ? _GEN_4136 : _GEN_4135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4138 = ~io_inputBit ? 1'h0 : _GEN_4137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4139 = i == 10'h282 ? _GEN_4138 : _GEN_4137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4140 = io_inputBit | _GEN_4139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4141 = i == 10'h282 ? _GEN_4140 : _GEN_4139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4142 = ~io_inputBit ? 1'h0 : _GEN_4141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4143 = i == 10'h283 ? _GEN_4142 : _GEN_4141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4144 = io_inputBit | _GEN_4143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4145 = i == 10'h283 ? _GEN_4144 : _GEN_4143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4146 = ~io_inputBit ? 1'h0 : _GEN_4145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4147 = i == 10'h284 ? _GEN_4146 : _GEN_4145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4148 = io_inputBit | _GEN_4147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4149 = i == 10'h284 ? _GEN_4148 : _GEN_4147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4150 = ~io_inputBit ? 1'h0 : _GEN_4149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4151 = i == 10'h285 ? _GEN_4150 : _GEN_4149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4152 = io_inputBit | _GEN_4151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4153 = i == 10'h285 ? _GEN_4152 : _GEN_4151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4154 = ~io_inputBit ? 1'h0 : _GEN_4153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4155 = i == 10'h286 ? _GEN_4154 : _GEN_4153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4156 = io_inputBit | _GEN_4155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4157 = i == 10'h286 ? _GEN_4156 : _GEN_4155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4158 = ~io_inputBit ? 1'h0 : _GEN_4157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4159 = i == 10'h287 ? _GEN_4158 : _GEN_4157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4160 = io_inputBit | _GEN_4159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4161 = i == 10'h287 ? _GEN_4160 : _GEN_4159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4162 = ~io_inputBit ? 1'h0 : _GEN_4161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4163 = i == 10'h288 ? _GEN_4162 : _GEN_4161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4164 = io_inputBit | _GEN_4163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4165 = i == 10'h288 ? _GEN_4164 : _GEN_4163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4166 = ~io_inputBit ? 1'h0 : _GEN_4165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4167 = i == 10'h289 ? _GEN_4166 : _GEN_4165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4168 = io_inputBit | _GEN_4167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4169 = i == 10'h289 ? _GEN_4168 : _GEN_4167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4170 = ~io_inputBit ? 1'h0 : _GEN_4169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4171 = i == 10'h28a ? _GEN_4170 : _GEN_4169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4172 = io_inputBit | _GEN_4171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4173 = i == 10'h28a ? _GEN_4172 : _GEN_4171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4174 = ~io_inputBit ? 1'h0 : _GEN_4173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4175 = i == 10'h28b ? _GEN_4174 : _GEN_4173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4176 = io_inputBit | _GEN_4175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4177 = i == 10'h28b ? _GEN_4176 : _GEN_4175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4178 = ~io_inputBit ? 1'h0 : _GEN_4177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4179 = i == 10'h28c ? _GEN_4178 : _GEN_4177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4180 = io_inputBit | _GEN_4179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4181 = i == 10'h28c ? _GEN_4180 : _GEN_4179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4182 = ~io_inputBit ? 1'h0 : _GEN_4181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4183 = i == 10'h28d ? _GEN_4182 : _GEN_4181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4184 = io_inputBit | _GEN_4183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4185 = i == 10'h28d ? _GEN_4184 : _GEN_4183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4186 = ~io_inputBit ? 1'h0 : _GEN_4185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4187 = i == 10'h28e ? _GEN_4186 : _GEN_4185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4188 = io_inputBit | _GEN_4187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4189 = i == 10'h28e ? _GEN_4188 : _GEN_4187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4190 = ~io_inputBit ? 1'h0 : _GEN_4189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4191 = i == 10'h28f ? _GEN_4190 : _GEN_4189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4192 = io_inputBit | _GEN_4191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4193 = i == 10'h28f ? _GEN_4192 : _GEN_4191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4194 = ~io_inputBit ? 1'h0 : _GEN_4193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4195 = i == 10'h290 ? _GEN_4194 : _GEN_4193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4196 = io_inputBit | _GEN_4195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4197 = i == 10'h290 ? _GEN_4196 : _GEN_4195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4198 = ~io_inputBit ? 1'h0 : _GEN_4197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4199 = i == 10'h291 ? _GEN_4198 : _GEN_4197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4200 = io_inputBit | _GEN_4199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4201 = i == 10'h291 ? _GEN_4200 : _GEN_4199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4202 = ~io_inputBit ? 1'h0 : _GEN_4201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4203 = i == 10'h292 ? _GEN_4202 : _GEN_4201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4204 = io_inputBit | _GEN_4203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4205 = i == 10'h292 ? _GEN_4204 : _GEN_4203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4206 = ~io_inputBit ? 1'h0 : _GEN_4205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4207 = i == 10'h293 ? _GEN_4206 : _GEN_4205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4208 = io_inputBit | _GEN_4207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4209 = i == 10'h293 ? _GEN_4208 : _GEN_4207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4210 = ~io_inputBit ? 1'h0 : _GEN_4209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4211 = i == 10'h294 ? _GEN_4210 : _GEN_4209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4212 = io_inputBit | _GEN_4211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4213 = i == 10'h294 ? _GEN_4212 : _GEN_4211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4214 = io_inputBit ? 1'h0 : _GEN_2807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4215 = i == 10'h0 ? _GEN_4214 : _GEN_2807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4216 = ~io_inputBit ? 1'h0 : _GEN_4215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4217 = i == 10'h1 ? _GEN_4216 : _GEN_4215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4218 = io_inputBit ? 1'h0 : _GEN_4217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4219 = i == 10'h4 ? _GEN_4218 : _GEN_4217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4220 = io_inputBit ? 1'h0 : _GEN_4219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4221 = i == 10'h9 ? _GEN_4220 : _GEN_4219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4222 = io_inputBit | _GEN_4221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4223 = i == 10'h27 ? _GEN_4222 : _GEN_4221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4224 = io_inputBit ? 1'h0 : _GEN_4223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4225 = i == 10'h28 ? _GEN_4224 : _GEN_4223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4226 = ~io_inputBit ? 1'h0 : _GEN_4225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4227 = i == 10'h4f ? _GEN_4226 : _GEN_4225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4228 = io_inputBit | _GEN_4227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4229 = i == 10'h4f ? _GEN_4228 : _GEN_4227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4230 = ~io_inputBit | _GEN_4229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4231 = i == 10'h51 ? _GEN_4230 : _GEN_4229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4232 = ~io_inputBit | _GEN_4231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4233 = i == 10'ha4 ? _GEN_4232 : _GEN_4231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4234 = io_inputBit ? 1'h0 : _GEN_4233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4235 = i == 10'h14a ? _GEN_4234 : _GEN_4233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4236 = ~io_inputBit | _GEN_4235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4237 = i == 10'h295 ? _GEN_4236 : _GEN_4235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4238 = io_inputBit ? 1'h0 : _GEN_4237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4239 = i == 10'h295 ? _GEN_4238 : _GEN_4237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4240 = io_inputBit ? 1'h0 : _GEN_2885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4241 = i == 10'h0 ? _GEN_4240 : _GEN_2885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4242 = ~io_inputBit ? 1'h0 : _GEN_4241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4243 = i == 10'h3 ? _GEN_4242 : _GEN_4241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4244 = io_inputBit ? 1'h0 : _GEN_4243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4245 = i == 10'h4 ? _GEN_4244 : _GEN_4243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4246 = ~io_inputBit ? 1'h0 : _GEN_4245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4247 = i == 10'h8 ? _GEN_4246 : _GEN_4245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4248 = io_inputBit ? 1'h0 : _GEN_4247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4249 = i == 10'h9 ? _GEN_4248 : _GEN_4247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4250 = ~io_inputBit ? 1'h0 : _GEN_4249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4251 = i == 10'h12 ? _GEN_4250 : _GEN_4249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4252 = io_inputBit | _GEN_4251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4253 = i == 10'h26 ? _GEN_4252 : _GEN_4251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4254 = io_inputBit ? 1'h0 : _GEN_4253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4255 = i == 10'h27 ? _GEN_4254 : _GEN_4253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4256 = io_inputBit ? 1'h0 : _GEN_4255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4257 = i == 10'h28 ? _GEN_4256 : _GEN_4255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4258 = ~io_inputBit ? 1'h0 : _GEN_4257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4259 = i == 10'h4d ? _GEN_4258 : _GEN_4257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4260 = io_inputBit | _GEN_4259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4261 = i == 10'h4d ? _GEN_4260 : _GEN_4259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4262 = ~io_inputBit | _GEN_4261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4263 = i == 10'h4f ? _GEN_4262 : _GEN_4261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4264 = io_inputBit ? 1'h0 : _GEN_4263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4265 = i == 10'h4f ? _GEN_4264 : _GEN_4263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4266 = ~io_inputBit ? 1'h0 : _GEN_4265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4267 = i == 10'h51 ? _GEN_4266 : _GEN_4265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4268 = ~io_inputBit | _GEN_4267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4269 = i == 10'ha4 ? _GEN_4268 : _GEN_4267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4270 = io_inputBit ? 1'h0 : _GEN_4269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4271 = i == 10'h14a ? _GEN_4270 : _GEN_4269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4272 = ~io_inputBit | _GEN_4271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4273 = i == 10'h295 ? _GEN_4272 : _GEN_4271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4274 = io_inputBit ? 1'h0 : _GEN_4273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4275 = i == 10'h295 ? _GEN_4274 : _GEN_4273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4276 = io_inputBit ? 1'h0 : _GEN_3005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4277 = i == 10'h0 ? _GEN_4276 : _GEN_3005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4278 = ~io_inputBit ? 1'h0 : _GEN_4277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4279 = i == 10'h3 ? _GEN_4278 : _GEN_4277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4280 = io_inputBit ? 1'h0 : _GEN_4279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4281 = i == 10'h4 ? _GEN_4280 : _GEN_4279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4282 = ~io_inputBit ? 1'h0 : _GEN_4281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4283 = i == 10'h8 ? _GEN_4282 : _GEN_4281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4284 = io_inputBit ? 1'h0 : _GEN_4283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4285 = i == 10'h9 ? _GEN_4284 : _GEN_4283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4286 = ~io_inputBit ? 1'h0 : _GEN_4285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4287 = i == 10'h25 ? _GEN_4286 : _GEN_4285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4288 = io_inputBit ? 1'h0 : _GEN_4287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4289 = i == 10'h28 ? _GEN_4288 : _GEN_4287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4290 = ~io_inputBit ? 1'h0 : _GEN_4289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4291 = i == 10'h4c ? _GEN_4290 : _GEN_4289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4292 = io_inputBit | _GEN_4291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4293 = i == 10'h4c ? _GEN_4292 : _GEN_4291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4294 = ~io_inputBit | _GEN_4293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4295 = i == 10'h4d ? _GEN_4294 : _GEN_4293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4296 = io_inputBit ? 1'h0 : _GEN_4295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4297 = i == 10'h4d ? _GEN_4296 : _GEN_4295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4298 = ~io_inputBit ? 1'h0 : _GEN_4297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4299 = i == 10'h4e ? _GEN_4298 : _GEN_4297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4300 = io_inputBit | _GEN_4299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4301 = i == 10'h4e ? _GEN_4300 : _GEN_4299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4302 = ~io_inputBit | _GEN_4301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4303 = i == 10'h4f ? _GEN_4302 : _GEN_4301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4304 = io_inputBit ? 1'h0 : _GEN_4303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4305 = i == 10'h4f ? _GEN_4304 : _GEN_4303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4306 = ~io_inputBit ? 1'h0 : _GEN_4305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4307 = i == 10'h50 ? _GEN_4306 : _GEN_4305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4308 = io_inputBit | _GEN_4307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4309 = i == 10'h50 ? _GEN_4308 : _GEN_4307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4310 = ~io_inputBit | _GEN_4309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4311 = i == 10'h51 ? _GEN_4310 : _GEN_4309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4312 = io_inputBit ? 1'h0 : _GEN_4311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4313 = i == 10'h51 ? _GEN_4312 : _GEN_4311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4314 = io_inputBit ? 1'h0 : _GEN_3195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4315 = i == 10'h0 ? _GEN_4314 : _GEN_3195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4316 = ~io_inputBit ? 1'h0 : _GEN_4315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4317 = i == 10'h3 ? _GEN_4316 : _GEN_4315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4318 = io_inputBit ? 1'h0 : _GEN_4317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4319 = i == 10'h4 ? _GEN_4318 : _GEN_4317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4320 = ~io_inputBit ? 1'h0 : _GEN_4319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4321 = i == 10'h8 ? _GEN_4320 : _GEN_4319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4322 = io_inputBit ? 1'h0 : _GEN_4321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4323 = i == 10'h9 ? _GEN_4322 : _GEN_4321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4324 = ~io_inputBit ? 1'h0 : _GEN_4323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4325 = i == 10'h25 ? _GEN_4324 : _GEN_4323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4326 = io_inputBit ? 1'h0 : _GEN_4325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4327 = i == 10'h28 ? _GEN_4326 : _GEN_4325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4328 = ~io_inputBit | _GEN_4327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4329 = i == 10'h4c ? _GEN_4328 : _GEN_4327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4330 = io_inputBit ? 1'h0 : _GEN_4329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4331 = i == 10'h4c ? _GEN_4330 : _GEN_4329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4332 = ~io_inputBit | _GEN_4331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4333 = i == 10'h4d ? _GEN_4332 : _GEN_4331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4334 = io_inputBit ? 1'h0 : _GEN_4333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4335 = i == 10'h4d ? _GEN_4334 : _GEN_4333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4336 = ~io_inputBit | _GEN_4335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4337 = i == 10'h4e ? _GEN_4336 : _GEN_4335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4338 = io_inputBit ? 1'h0 : _GEN_4337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4339 = i == 10'h4e ? _GEN_4338 : _GEN_4337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4340 = ~io_inputBit | _GEN_4339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4341 = i == 10'h4f ? _GEN_4340 : _GEN_4339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4342 = io_inputBit ? 1'h0 : _GEN_4341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4343 = i == 10'h4f ? _GEN_4342 : _GEN_4341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4344 = ~io_inputBit | _GEN_4343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4345 = i == 10'h50 ? _GEN_4344 : _GEN_4343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4346 = io_inputBit ? 1'h0 : _GEN_4345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4347 = i == 10'h50 ? _GEN_4346 : _GEN_4345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4348 = ~io_inputBit | _GEN_4347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4349 = i == 10'h51 ? _GEN_4348 : _GEN_4347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4350 = io_inputBit ? 1'h0 : _GEN_4349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4351 = i == 10'h51 ? _GEN_4350 : _GEN_4349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4352 = io_inputBit ? 1'h0 : _GEN_3467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4353 = i == 10'h0 ? _GEN_4352 : _GEN_3467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4354 = ~io_inputBit ? 1'h0 : _GEN_4353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4355 = i == 10'h3 ? _GEN_4354 : _GEN_4353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4356 = io_inputBit ? 1'h0 : _GEN_4355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4357 = i == 10'h4 ? _GEN_4356 : _GEN_4355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4358 = ~io_inputBit ? 1'h0 : _GEN_4357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4359 = i == 10'h8 ? _GEN_4358 : _GEN_4357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4360 = io_inputBit ? 1'h0 : _GEN_4359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4361 = i == 10'h9 ? _GEN_4360 : _GEN_4359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4362 = io_inputBit ? 1'h0 : _GEN_4361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4363 = i == 10'h28 ? _GEN_4362 : _GEN_4361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4364 = ~io_inputBit ? 1'h0 : _GEN_4363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4365 = i == 10'h4b ? _GEN_4364 : _GEN_4363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4366 = ~io_inputBit ? 1'h0 : _GEN_4365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4367 = i == 10'h98 ? _GEN_4366 : _GEN_4365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4368 = io_inputBit | _GEN_4367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4369 = i == 10'h98 ? _GEN_4368 : _GEN_4367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4370 = ~io_inputBit ? 1'h0 : _GEN_4369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4371 = i == 10'h99 ? _GEN_4370 : _GEN_4369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4372 = io_inputBit | _GEN_4371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4373 = i == 10'h99 ? _GEN_4372 : _GEN_4371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4374 = ~io_inputBit ? 1'h0 : _GEN_4373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4375 = i == 10'h9a ? _GEN_4374 : _GEN_4373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4376 = io_inputBit | _GEN_4375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4377 = i == 10'h9a ? _GEN_4376 : _GEN_4375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4378 = ~io_inputBit ? 1'h0 : _GEN_4377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4379 = i == 10'h9b ? _GEN_4378 : _GEN_4377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4380 = io_inputBit | _GEN_4379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4381 = i == 10'h9b ? _GEN_4380 : _GEN_4379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4382 = ~io_inputBit ? 1'h0 : _GEN_4381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4383 = i == 10'h9c ? _GEN_4382 : _GEN_4381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4384 = io_inputBit | _GEN_4383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4385 = i == 10'h9c ? _GEN_4384 : _GEN_4383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4386 = ~io_inputBit ? 1'h0 : _GEN_4385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4387 = i == 10'h9d ? _GEN_4386 : _GEN_4385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4388 = io_inputBit | _GEN_4387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4389 = i == 10'h9d ? _GEN_4388 : _GEN_4387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4390 = ~io_inputBit ? 1'h0 : _GEN_4389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4391 = i == 10'h9e ? _GEN_4390 : _GEN_4389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4392 = io_inputBit | _GEN_4391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4393 = i == 10'h9e ? _GEN_4392 : _GEN_4391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4394 = ~io_inputBit ? 1'h0 : _GEN_4393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4395 = i == 10'h9f ? _GEN_4394 : _GEN_4393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4396 = io_inputBit | _GEN_4395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4397 = i == 10'h9f ? _GEN_4396 : _GEN_4395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4398 = ~io_inputBit ? 1'h0 : _GEN_4397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4399 = i == 10'ha0 ? _GEN_4398 : _GEN_4397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4400 = io_inputBit | _GEN_4399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4401 = i == 10'ha0 ? _GEN_4400 : _GEN_4399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4402 = ~io_inputBit ? 1'h0 : _GEN_4401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4403 = i == 10'ha1 ? _GEN_4402 : _GEN_4401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4404 = io_inputBit | _GEN_4403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4405 = i == 10'ha1 ? _GEN_4404 : _GEN_4403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4406 = ~io_inputBit ? 1'h0 : _GEN_4405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4407 = i == 10'ha2 ? _GEN_4406 : _GEN_4405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4408 = io_inputBit | _GEN_4407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4409 = i == 10'ha2 ? _GEN_4408 : _GEN_4407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4410 = ~io_inputBit ? 1'h0 : _GEN_4409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4411 = i == 10'ha3 ? _GEN_4410 : _GEN_4409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4412 = io_inputBit | _GEN_4411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4413 = i == 10'ha3 ? _GEN_4412 : _GEN_4411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4414 = ~io_inputBit ? 1'h0 : _GEN_4413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4415 = i == 10'ha4 ? _GEN_4414 : _GEN_4413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4416 = io_inputBit ? 1'h0 : _GEN_4415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4417 = i == 10'h14a ? _GEN_4416 : _GEN_4415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4418 = ~io_inputBit | _GEN_4417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4419 = i == 10'h295 ? _GEN_4418 : _GEN_4417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4420 = io_inputBit ? 1'h0 : _GEN_4419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4421 = i == 10'h295 ? _GEN_4420 : _GEN_4419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4422 = io_inputBit ? 1'h0 : _GEN_3789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4423 = i == 10'h0 ? _GEN_4422 : _GEN_3789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4424 = ~io_inputBit ? 1'h0 : _GEN_4423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4425 = i == 10'h3 ? _GEN_4424 : _GEN_4423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4426 = io_inputBit ? 1'h0 : _GEN_4425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4427 = i == 10'h4 ? _GEN_4426 : _GEN_4425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4428 = ~io_inputBit ? 1'h0 : _GEN_4427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4429 = i == 10'h8 ? _GEN_4428 : _GEN_4427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4430 = io_inputBit ? 1'h0 : _GEN_4429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4431 = i == 10'h9 ? _GEN_4430 : _GEN_4429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4432 = io_inputBit ? 1'h0 : _GEN_4431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4433 = i == 10'h28 ? _GEN_4432 : _GEN_4431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4434 = ~io_inputBit ? 1'h0 : _GEN_4433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4435 = i == 10'h4b ? _GEN_4434 : _GEN_4433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4436 = io_inputBit ? 1'h0 : _GEN_4435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4437 = i == 10'ha4 ? _GEN_4436 : _GEN_4435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4438 = ~io_inputBit ? 1'h0 : _GEN_4437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4439 = i == 10'h131 ? _GEN_4438 : _GEN_4437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4440 = io_inputBit | _GEN_4439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4441 = i == 10'h131 ? _GEN_4440 : _GEN_4439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4442 = ~io_inputBit ? 1'h0 : _GEN_4441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4443 = i == 10'h132 ? _GEN_4442 : _GEN_4441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4444 = io_inputBit | _GEN_4443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4445 = i == 10'h132 ? _GEN_4444 : _GEN_4443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4446 = ~io_inputBit ? 1'h0 : _GEN_4445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4447 = i == 10'h133 ? _GEN_4446 : _GEN_4445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4448 = io_inputBit | _GEN_4447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4449 = i == 10'h133 ? _GEN_4448 : _GEN_4447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4450 = ~io_inputBit ? 1'h0 : _GEN_4449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4451 = i == 10'h134 ? _GEN_4450 : _GEN_4449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4452 = io_inputBit | _GEN_4451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4453 = i == 10'h134 ? _GEN_4452 : _GEN_4451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4454 = ~io_inputBit ? 1'h0 : _GEN_4453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4455 = i == 10'h135 ? _GEN_4454 : _GEN_4453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4456 = io_inputBit | _GEN_4455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4457 = i == 10'h135 ? _GEN_4456 : _GEN_4455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4458 = ~io_inputBit ? 1'h0 : _GEN_4457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4459 = i == 10'h136 ? _GEN_4458 : _GEN_4457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4460 = io_inputBit | _GEN_4459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4461 = i == 10'h136 ? _GEN_4460 : _GEN_4459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4462 = ~io_inputBit ? 1'h0 : _GEN_4461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4463 = i == 10'h137 ? _GEN_4462 : _GEN_4461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4464 = io_inputBit | _GEN_4463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4465 = i == 10'h137 ? _GEN_4464 : _GEN_4463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4466 = ~io_inputBit ? 1'h0 : _GEN_4465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4467 = i == 10'h138 ? _GEN_4466 : _GEN_4465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4468 = io_inputBit | _GEN_4467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4469 = i == 10'h138 ? _GEN_4468 : _GEN_4467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4470 = ~io_inputBit ? 1'h0 : _GEN_4469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4471 = i == 10'h139 ? _GEN_4470 : _GEN_4469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4472 = io_inputBit | _GEN_4471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4473 = i == 10'h139 ? _GEN_4472 : _GEN_4471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4474 = ~io_inputBit ? 1'h0 : _GEN_4473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4475 = i == 10'h13a ? _GEN_4474 : _GEN_4473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4476 = io_inputBit | _GEN_4475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4477 = i == 10'h13a ? _GEN_4476 : _GEN_4475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4478 = ~io_inputBit ? 1'h0 : _GEN_4477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4479 = i == 10'h13b ? _GEN_4478 : _GEN_4477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4480 = io_inputBit | _GEN_4479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4481 = i == 10'h13b ? _GEN_4480 : _GEN_4479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4482 = ~io_inputBit ? 1'h0 : _GEN_4481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4483 = i == 10'h13c ? _GEN_4482 : _GEN_4481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4484 = io_inputBit | _GEN_4483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4485 = i == 10'h13c ? _GEN_4484 : _GEN_4483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4486 = ~io_inputBit ? 1'h0 : _GEN_4485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4487 = i == 10'h13d ? _GEN_4486 : _GEN_4485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4488 = io_inputBit | _GEN_4487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4489 = i == 10'h13d ? _GEN_4488 : _GEN_4487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4490 = ~io_inputBit ? 1'h0 : _GEN_4489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4491 = i == 10'h13e ? _GEN_4490 : _GEN_4489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4492 = io_inputBit | _GEN_4491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4493 = i == 10'h13e ? _GEN_4492 : _GEN_4491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4494 = ~io_inputBit ? 1'h0 : _GEN_4493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4495 = i == 10'h13f ? _GEN_4494 : _GEN_4493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4496 = io_inputBit | _GEN_4495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4497 = i == 10'h13f ? _GEN_4496 : _GEN_4495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4498 = ~io_inputBit ? 1'h0 : _GEN_4497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4499 = i == 10'h140 ? _GEN_4498 : _GEN_4497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4500 = io_inputBit | _GEN_4499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4501 = i == 10'h140 ? _GEN_4500 : _GEN_4499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4502 = ~io_inputBit ? 1'h0 : _GEN_4501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4503 = i == 10'h141 ? _GEN_4502 : _GEN_4501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4504 = io_inputBit | _GEN_4503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4505 = i == 10'h141 ? _GEN_4504 : _GEN_4503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4506 = ~io_inputBit ? 1'h0 : _GEN_4505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4507 = i == 10'h142 ? _GEN_4506 : _GEN_4505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4508 = io_inputBit | _GEN_4507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4509 = i == 10'h142 ? _GEN_4508 : _GEN_4507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4510 = ~io_inputBit ? 1'h0 : _GEN_4509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4511 = i == 10'h143 ? _GEN_4510 : _GEN_4509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4512 = io_inputBit | _GEN_4511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4513 = i == 10'h143 ? _GEN_4512 : _GEN_4511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4514 = ~io_inputBit ? 1'h0 : _GEN_4513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4515 = i == 10'h144 ? _GEN_4514 : _GEN_4513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4516 = io_inputBit | _GEN_4515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4517 = i == 10'h144 ? _GEN_4516 : _GEN_4515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4518 = ~io_inputBit ? 1'h0 : _GEN_4517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4519 = i == 10'h145 ? _GEN_4518 : _GEN_4517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4520 = io_inputBit | _GEN_4519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4521 = i == 10'h145 ? _GEN_4520 : _GEN_4519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4522 = ~io_inputBit ? 1'h0 : _GEN_4521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4523 = i == 10'h146 ? _GEN_4522 : _GEN_4521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4524 = io_inputBit | _GEN_4523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4525 = i == 10'h146 ? _GEN_4524 : _GEN_4523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4526 = ~io_inputBit ? 1'h0 : _GEN_4525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4527 = i == 10'h147 ? _GEN_4526 : _GEN_4525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4528 = io_inputBit | _GEN_4527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4529 = i == 10'h147 ? _GEN_4528 : _GEN_4527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4530 = ~io_inputBit ? 1'h0 : _GEN_4529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4531 = i == 10'h148 ? _GEN_4530 : _GEN_4529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4532 = io_inputBit | _GEN_4531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4533 = i == 10'h148 ? _GEN_4532 : _GEN_4531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4534 = ~io_inputBit ? 1'h0 : _GEN_4533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4535 = i == 10'h149 ? _GEN_4534 : _GEN_4533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4536 = io_inputBit | _GEN_4535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4537 = i == 10'h149 ? _GEN_4536 : _GEN_4535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4538 = io_inputBit ? 1'h0 : _GEN_4213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4539 = i == 10'h0 ? _GEN_4538 : _GEN_4213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4540 = ~io_inputBit ? 1'h0 : _GEN_4539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4541 = i == 10'h3 ? _GEN_4540 : _GEN_4539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4542 = io_inputBit ? 1'h0 : _GEN_4541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4543 = i == 10'h4 ? _GEN_4542 : _GEN_4541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4544 = ~io_inputBit ? 1'h0 : _GEN_4543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4545 = i == 10'h8 ? _GEN_4544 : _GEN_4543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4546 = io_inputBit ? 1'h0 : _GEN_4545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4547 = i == 10'h9 ? _GEN_4546 : _GEN_4545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4548 = io_inputBit ? 1'h0 : _GEN_4547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4549 = i == 10'h28 ? _GEN_4548 : _GEN_4547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4550 = ~io_inputBit ? 1'h0 : _GEN_4549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4551 = i == 10'h4b ? _GEN_4550 : _GEN_4549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4552 = io_inputBit ? 1'h0 : _GEN_4551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4553 = i == 10'ha4 ? _GEN_4552 : _GEN_4551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4554 = ~io_inputBit ? 1'h0 : _GEN_4553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4555 = i == 10'h263 ? _GEN_4554 : _GEN_4553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4556 = io_inputBit | _GEN_4555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4557 = i == 10'h263 ? _GEN_4556 : _GEN_4555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4558 = ~io_inputBit ? 1'h0 : _GEN_4557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4559 = i == 10'h264 ? _GEN_4558 : _GEN_4557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4560 = io_inputBit | _GEN_4559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4561 = i == 10'h264 ? _GEN_4560 : _GEN_4559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4562 = ~io_inputBit ? 1'h0 : _GEN_4561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4563 = i == 10'h265 ? _GEN_4562 : _GEN_4561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4564 = io_inputBit | _GEN_4563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4565 = i == 10'h265 ? _GEN_4564 : _GEN_4563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4566 = ~io_inputBit ? 1'h0 : _GEN_4565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4567 = i == 10'h266 ? _GEN_4566 : _GEN_4565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4568 = io_inputBit | _GEN_4567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4569 = i == 10'h266 ? _GEN_4568 : _GEN_4567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4570 = ~io_inputBit ? 1'h0 : _GEN_4569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4571 = i == 10'h267 ? _GEN_4570 : _GEN_4569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4572 = io_inputBit | _GEN_4571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4573 = i == 10'h267 ? _GEN_4572 : _GEN_4571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4574 = ~io_inputBit ? 1'h0 : _GEN_4573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4575 = i == 10'h268 ? _GEN_4574 : _GEN_4573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4576 = io_inputBit | _GEN_4575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4577 = i == 10'h268 ? _GEN_4576 : _GEN_4575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4578 = ~io_inputBit ? 1'h0 : _GEN_4577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4579 = i == 10'h269 ? _GEN_4578 : _GEN_4577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4580 = io_inputBit | _GEN_4579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4581 = i == 10'h269 ? _GEN_4580 : _GEN_4579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4582 = ~io_inputBit ? 1'h0 : _GEN_4581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4583 = i == 10'h26a ? _GEN_4582 : _GEN_4581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4584 = io_inputBit | _GEN_4583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4585 = i == 10'h26a ? _GEN_4584 : _GEN_4583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4586 = ~io_inputBit ? 1'h0 : _GEN_4585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4587 = i == 10'h26b ? _GEN_4586 : _GEN_4585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4588 = io_inputBit | _GEN_4587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4589 = i == 10'h26b ? _GEN_4588 : _GEN_4587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4590 = ~io_inputBit ? 1'h0 : _GEN_4589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4591 = i == 10'h26c ? _GEN_4590 : _GEN_4589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4592 = io_inputBit | _GEN_4591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4593 = i == 10'h26c ? _GEN_4592 : _GEN_4591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4594 = ~io_inputBit ? 1'h0 : _GEN_4593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4595 = i == 10'h26d ? _GEN_4594 : _GEN_4593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4596 = io_inputBit | _GEN_4595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4597 = i == 10'h26d ? _GEN_4596 : _GEN_4595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4598 = ~io_inputBit ? 1'h0 : _GEN_4597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4599 = i == 10'h26e ? _GEN_4598 : _GEN_4597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4600 = io_inputBit | _GEN_4599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4601 = i == 10'h26e ? _GEN_4600 : _GEN_4599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4602 = ~io_inputBit ? 1'h0 : _GEN_4601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4603 = i == 10'h26f ? _GEN_4602 : _GEN_4601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4604 = io_inputBit | _GEN_4603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4605 = i == 10'h26f ? _GEN_4604 : _GEN_4603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4606 = ~io_inputBit ? 1'h0 : _GEN_4605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4607 = i == 10'h270 ? _GEN_4606 : _GEN_4605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4608 = io_inputBit | _GEN_4607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4609 = i == 10'h270 ? _GEN_4608 : _GEN_4607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4610 = ~io_inputBit ? 1'h0 : _GEN_4609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4611 = i == 10'h271 ? _GEN_4610 : _GEN_4609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4612 = io_inputBit | _GEN_4611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4613 = i == 10'h271 ? _GEN_4612 : _GEN_4611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4614 = ~io_inputBit ? 1'h0 : _GEN_4613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4615 = i == 10'h272 ? _GEN_4614 : _GEN_4613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4616 = io_inputBit | _GEN_4615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4617 = i == 10'h272 ? _GEN_4616 : _GEN_4615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4618 = ~io_inputBit ? 1'h0 : _GEN_4617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4619 = i == 10'h273 ? _GEN_4618 : _GEN_4617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4620 = io_inputBit | _GEN_4619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4621 = i == 10'h273 ? _GEN_4620 : _GEN_4619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4622 = ~io_inputBit ? 1'h0 : _GEN_4621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4623 = i == 10'h274 ? _GEN_4622 : _GEN_4621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4624 = io_inputBit | _GEN_4623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4625 = i == 10'h274 ? _GEN_4624 : _GEN_4623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4626 = ~io_inputBit ? 1'h0 : _GEN_4625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4627 = i == 10'h275 ? _GEN_4626 : _GEN_4625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4628 = io_inputBit | _GEN_4627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4629 = i == 10'h275 ? _GEN_4628 : _GEN_4627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4630 = ~io_inputBit ? 1'h0 : _GEN_4629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4631 = i == 10'h276 ? _GEN_4630 : _GEN_4629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4632 = io_inputBit | _GEN_4631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4633 = i == 10'h276 ? _GEN_4632 : _GEN_4631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4634 = ~io_inputBit ? 1'h0 : _GEN_4633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4635 = i == 10'h277 ? _GEN_4634 : _GEN_4633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4636 = io_inputBit | _GEN_4635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4637 = i == 10'h277 ? _GEN_4636 : _GEN_4635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4638 = ~io_inputBit ? 1'h0 : _GEN_4637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4639 = i == 10'h278 ? _GEN_4638 : _GEN_4637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4640 = io_inputBit | _GEN_4639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4641 = i == 10'h278 ? _GEN_4640 : _GEN_4639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4642 = ~io_inputBit ? 1'h0 : _GEN_4641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4643 = i == 10'h279 ? _GEN_4642 : _GEN_4641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4644 = io_inputBit | _GEN_4643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4645 = i == 10'h279 ? _GEN_4644 : _GEN_4643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4646 = ~io_inputBit ? 1'h0 : _GEN_4645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4647 = i == 10'h27a ? _GEN_4646 : _GEN_4645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4648 = io_inputBit | _GEN_4647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4649 = i == 10'h27a ? _GEN_4648 : _GEN_4647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4650 = ~io_inputBit ? 1'h0 : _GEN_4649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4651 = i == 10'h27b ? _GEN_4650 : _GEN_4649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4652 = io_inputBit | _GEN_4651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4653 = i == 10'h27b ? _GEN_4652 : _GEN_4651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4654 = ~io_inputBit ? 1'h0 : _GEN_4653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4655 = i == 10'h27c ? _GEN_4654 : _GEN_4653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4656 = io_inputBit | _GEN_4655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4657 = i == 10'h27c ? _GEN_4656 : _GEN_4655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4658 = ~io_inputBit ? 1'h0 : _GEN_4657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4659 = i == 10'h27d ? _GEN_4658 : _GEN_4657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4660 = io_inputBit | _GEN_4659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4661 = i == 10'h27d ? _GEN_4660 : _GEN_4659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4662 = ~io_inputBit ? 1'h0 : _GEN_4661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4663 = i == 10'h27e ? _GEN_4662 : _GEN_4661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4664 = io_inputBit | _GEN_4663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4665 = i == 10'h27e ? _GEN_4664 : _GEN_4663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4666 = ~io_inputBit ? 1'h0 : _GEN_4665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4667 = i == 10'h27f ? _GEN_4666 : _GEN_4665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4668 = io_inputBit | _GEN_4667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4669 = i == 10'h27f ? _GEN_4668 : _GEN_4667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4670 = ~io_inputBit ? 1'h0 : _GEN_4669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4671 = i == 10'h280 ? _GEN_4670 : _GEN_4669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4672 = io_inputBit | _GEN_4671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4673 = i == 10'h280 ? _GEN_4672 : _GEN_4671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4674 = ~io_inputBit ? 1'h0 : _GEN_4673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4675 = i == 10'h281 ? _GEN_4674 : _GEN_4673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4676 = io_inputBit | _GEN_4675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4677 = i == 10'h281 ? _GEN_4676 : _GEN_4675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4678 = ~io_inputBit ? 1'h0 : _GEN_4677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4679 = i == 10'h282 ? _GEN_4678 : _GEN_4677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4680 = io_inputBit | _GEN_4679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4681 = i == 10'h282 ? _GEN_4680 : _GEN_4679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4682 = ~io_inputBit ? 1'h0 : _GEN_4681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4683 = i == 10'h283 ? _GEN_4682 : _GEN_4681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4684 = io_inputBit | _GEN_4683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4685 = i == 10'h283 ? _GEN_4684 : _GEN_4683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4686 = ~io_inputBit ? 1'h0 : _GEN_4685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4687 = i == 10'h284 ? _GEN_4686 : _GEN_4685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4688 = io_inputBit | _GEN_4687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4689 = i == 10'h284 ? _GEN_4688 : _GEN_4687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4690 = ~io_inputBit ? 1'h0 : _GEN_4689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4691 = i == 10'h285 ? _GEN_4690 : _GEN_4689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4692 = io_inputBit | _GEN_4691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4693 = i == 10'h285 ? _GEN_4692 : _GEN_4691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4694 = ~io_inputBit ? 1'h0 : _GEN_4693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4695 = i == 10'h286 ? _GEN_4694 : _GEN_4693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4696 = io_inputBit | _GEN_4695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4697 = i == 10'h286 ? _GEN_4696 : _GEN_4695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4698 = ~io_inputBit ? 1'h0 : _GEN_4697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4699 = i == 10'h287 ? _GEN_4698 : _GEN_4697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4700 = io_inputBit | _GEN_4699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4701 = i == 10'h287 ? _GEN_4700 : _GEN_4699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4702 = ~io_inputBit ? 1'h0 : _GEN_4701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4703 = i == 10'h288 ? _GEN_4702 : _GEN_4701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4704 = io_inputBit | _GEN_4703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4705 = i == 10'h288 ? _GEN_4704 : _GEN_4703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4706 = ~io_inputBit ? 1'h0 : _GEN_4705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4707 = i == 10'h289 ? _GEN_4706 : _GEN_4705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4708 = io_inputBit | _GEN_4707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4709 = i == 10'h289 ? _GEN_4708 : _GEN_4707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4710 = ~io_inputBit ? 1'h0 : _GEN_4709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4711 = i == 10'h28a ? _GEN_4710 : _GEN_4709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4712 = io_inputBit | _GEN_4711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4713 = i == 10'h28a ? _GEN_4712 : _GEN_4711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4714 = ~io_inputBit ? 1'h0 : _GEN_4713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4715 = i == 10'h28b ? _GEN_4714 : _GEN_4713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4716 = io_inputBit | _GEN_4715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4717 = i == 10'h28b ? _GEN_4716 : _GEN_4715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4718 = ~io_inputBit ? 1'h0 : _GEN_4717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4719 = i == 10'h28c ? _GEN_4718 : _GEN_4717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4720 = io_inputBit | _GEN_4719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4721 = i == 10'h28c ? _GEN_4720 : _GEN_4719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4722 = ~io_inputBit ? 1'h0 : _GEN_4721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4723 = i == 10'h28d ? _GEN_4722 : _GEN_4721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4724 = io_inputBit | _GEN_4723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4725 = i == 10'h28d ? _GEN_4724 : _GEN_4723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4726 = ~io_inputBit ? 1'h0 : _GEN_4725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4727 = i == 10'h28e ? _GEN_4726 : _GEN_4725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4728 = io_inputBit | _GEN_4727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4729 = i == 10'h28e ? _GEN_4728 : _GEN_4727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4730 = ~io_inputBit ? 1'h0 : _GEN_4729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4731 = i == 10'h28f ? _GEN_4730 : _GEN_4729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4732 = io_inputBit | _GEN_4731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4733 = i == 10'h28f ? _GEN_4732 : _GEN_4731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4734 = ~io_inputBit ? 1'h0 : _GEN_4733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4735 = i == 10'h290 ? _GEN_4734 : _GEN_4733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4736 = io_inputBit | _GEN_4735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4737 = i == 10'h290 ? _GEN_4736 : _GEN_4735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4738 = ~io_inputBit ? 1'h0 : _GEN_4737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4739 = i == 10'h291 ? _GEN_4738 : _GEN_4737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4740 = io_inputBit | _GEN_4739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4741 = i == 10'h291 ? _GEN_4740 : _GEN_4739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4742 = ~io_inputBit ? 1'h0 : _GEN_4741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4743 = i == 10'h292 ? _GEN_4742 : _GEN_4741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4744 = io_inputBit | _GEN_4743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4745 = i == 10'h292 ? _GEN_4744 : _GEN_4743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4746 = ~io_inputBit ? 1'h0 : _GEN_4745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4747 = i == 10'h293 ? _GEN_4746 : _GEN_4745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4748 = io_inputBit | _GEN_4747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4749 = i == 10'h293 ? _GEN_4748 : _GEN_4747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4750 = ~io_inputBit ? 1'h0 : _GEN_4749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4751 = i == 10'h294 ? _GEN_4750 : _GEN_4749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4752 = io_inputBit | _GEN_4751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4753 = i == 10'h294 ? _GEN_4752 : _GEN_4751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4754 = io_inputBit ? 1'h0 : _GEN_4239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4755 = i == 10'h0 ? _GEN_4754 : _GEN_4239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4756 = ~io_inputBit ? 1'h0 : _GEN_4755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4757 = i == 10'h1 ? _GEN_4756 : _GEN_4755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4758 = ~io_inputBit ? 1'h0 : _GEN_4757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4759 = i == 10'h4 ? _GEN_4758 : _GEN_4757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4760 = io_inputBit | _GEN_4759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4761 = i == 10'h15 ? _GEN_4760 : _GEN_4759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4762 = ~io_inputBit | _GEN_4761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4763 = i == 10'h16 ? _GEN_4762 : _GEN_4761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4764 = ~io_inputBit ? 1'h0 : _GEN_4763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4765 = i == 10'h2b ? _GEN_4764 : _GEN_4763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4766 = io_inputBit ? 1'h0 : _GEN_4765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4767 = i == 10'h2e ? _GEN_4766 : _GEN_4765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4768 = ~io_inputBit ? 1'h0 : _GEN_4767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4769 = i == 10'h58 ? _GEN_4768 : _GEN_4767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4770 = io_inputBit ? 1'h0 : _GEN_4769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4771 = i == 10'h5d ? _GEN_4770 : _GEN_4769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4772 = ~io_inputBit ? 1'h0 : _GEN_4771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4773 = i == 10'hb2 ? _GEN_4772 : _GEN_4771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4774 = ~io_inputBit | _GEN_4773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4775 = i == 10'hbb ? _GEN_4774 : _GEN_4773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4776 = ~io_inputBit ? 1'h0 : _GEN_4775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4777 = i == 10'h166 ? _GEN_4776 : _GEN_4775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4778 = io_inputBit | _GEN_4777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4779 = i == 10'h166 ? _GEN_4778 : _GEN_4777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4780 = ~io_inputBit | _GEN_4779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4781 = i == 10'h178 ? _GEN_4780 : _GEN_4779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4782 = ~io_inputBit | _GEN_4781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4783 = i == 10'h2f2 ? _GEN_4782 : _GEN_4781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4784 = io_inputBit ? 1'h0 : _GEN_4783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4785 = i == 10'h2f2 ? _GEN_4784 : _GEN_4783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4786 = ~io_inputBit ? 1'h0 : _GEN_4275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4787 = i == 10'h1 ? _GEN_4786 : _GEN_4275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4788 = io_inputBit ? 1'h0 : _GEN_4787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4789 = i == 10'h2 ? _GEN_4788 : _GEN_4787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4790 = io_inputBit ? 1'h0 : _GEN_4789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4791 = i == 10'h5 ? _GEN_4790 : _GEN_4789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4792 = ~io_inputBit ? 1'h0 : _GEN_4791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4793 = i == 10'h9 ? _GEN_4792 : _GEN_4791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4794 = io_inputBit ? 1'h0 : _GEN_4793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4795 = i == 10'hb ? _GEN_4794 : _GEN_4793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4796 = ~io_inputBit ? 1'h0 : _GEN_4795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4797 = i == 10'h14 ? _GEN_4796 : _GEN_4795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4798 = io_inputBit ? 1'h0 : _GEN_4797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4799 = i == 10'h17 ? _GEN_4798 : _GEN_4797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4800 = ~io_inputBit ? 1'h0 : _GEN_4799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4801 = i == 10'h2a ? _GEN_4800 : _GEN_4799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4802 = ~io_inputBit | _GEN_4801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4803 = i == 10'h2b ? _GEN_4802 : _GEN_4801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4804 = ~io_inputBit ? 1'h0 : _GEN_4803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4805 = i == 10'h2c ? _GEN_4804 : _GEN_4803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4806 = io_inputBit ? 1'h0 : _GEN_4805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4807 = i == 10'h2d ? _GEN_4806 : _GEN_4805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4808 = io_inputBit | _GEN_4807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4809 = i == 10'h2e ? _GEN_4808 : _GEN_4807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4810 = io_inputBit ? 1'h0 : _GEN_4809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4811 = i == 10'h2f ? _GEN_4810 : _GEN_4809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4812 = ~io_inputBit ? 1'h0 : _GEN_4811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4813 = i == 10'h56 ? _GEN_4812 : _GEN_4811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4814 = ~io_inputBit | _GEN_4813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4815 = i == 10'h58 ? _GEN_4814 : _GEN_4813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4816 = ~io_inputBit ? 1'h0 : _GEN_4815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4817 = i == 10'h5a ? _GEN_4816 : _GEN_4815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4818 = io_inputBit ? 1'h0 : _GEN_4817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4819 = i == 10'h5b ? _GEN_4818 : _GEN_4817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4820 = io_inputBit | _GEN_4819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4821 = i == 10'h5d ? _GEN_4820 : _GEN_4819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4822 = io_inputBit ? 1'h0 : _GEN_4821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4823 = i == 10'h5f ? _GEN_4822 : _GEN_4821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4824 = ~io_inputBit ? 1'h0 : _GEN_4823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4825 = i == 10'hae ? _GEN_4824 : _GEN_4823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4826 = ~io_inputBit | _GEN_4825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4827 = i == 10'hb2 ? _GEN_4826 : _GEN_4825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4828 = ~io_inputBit ? 1'h0 : _GEN_4827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4829 = i == 10'hb6 ? _GEN_4828 : _GEN_4827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4830 = ~io_inputBit | _GEN_4829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4831 = i == 10'hb7 ? _GEN_4830 : _GEN_4829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4832 = ~io_inputBit ? 1'h0 : _GEN_4831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4833 = i == 10'hbb ? _GEN_4832 : _GEN_4831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4834 = ~io_inputBit | _GEN_4833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4835 = i == 10'hbf ? _GEN_4834 : _GEN_4833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4836 = ~io_inputBit ? 1'h0 : _GEN_4835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4837 = i == 10'h15e ? _GEN_4836 : _GEN_4835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4838 = io_inputBit | _GEN_4837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4839 = i == 10'h15e ? _GEN_4838 : _GEN_4837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4840 = ~io_inputBit | _GEN_4839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4841 = i == 10'h166 ? _GEN_4840 : _GEN_4839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4842 = io_inputBit ? 1'h0 : _GEN_4841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4843 = i == 10'h166 ? _GEN_4842 : _GEN_4841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4844 = ~io_inputBit ? 1'h0 : _GEN_4843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4845 = i == 10'h16e ? _GEN_4844 : _GEN_4843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4846 = io_inputBit | _GEN_4845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4847 = i == 10'h16e ? _GEN_4846 : _GEN_4845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4848 = ~io_inputBit | _GEN_4847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4849 = i == 10'h170 ? _GEN_4848 : _GEN_4847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4850 = ~io_inputBit ? 1'h0 : _GEN_4849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4851 = i == 10'h178 ? _GEN_4850 : _GEN_4849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4852 = ~io_inputBit | _GEN_4851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4853 = i == 10'h180 ? _GEN_4852 : _GEN_4851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4854 = ~io_inputBit | _GEN_4853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4855 = i == 10'h2e2 ? _GEN_4854 : _GEN_4853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4856 = io_inputBit ? 1'h0 : _GEN_4855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4857 = i == 10'h2e2 ? _GEN_4856 : _GEN_4855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4858 = ~io_inputBit ? 1'h0 : _GEN_4857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4859 = i == 10'h2f2 ? _GEN_4858 : _GEN_4857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4860 = io_inputBit | _GEN_4859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4861 = i == 10'h2f2 ? _GEN_4860 : _GEN_4859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4862 = ~io_inputBit | _GEN_4861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4863 = i == 10'h302 ? _GEN_4862 : _GEN_4861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4864 = io_inputBit ? 1'h0 : _GEN_4863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4865 = i == 10'h302 ? _GEN_4864 : _GEN_4863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4866 = ~io_inputBit ? 1'h0 : _GEN_4313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4867 = i == 10'h1 ? _GEN_4866 : _GEN_4313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4868 = io_inputBit ? 1'h0 : _GEN_4867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4869 = i == 10'h2 ? _GEN_4868 : _GEN_4867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4870 = io_inputBit ? 1'h0 : _GEN_4869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4871 = i == 10'h5 ? _GEN_4870 : _GEN_4869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4872 = ~io_inputBit ? 1'h0 : _GEN_4871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4873 = i == 10'h9 ? _GEN_4872 : _GEN_4871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4874 = io_inputBit ? 1'h0 : _GEN_4873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4875 = i == 10'hb ? _GEN_4874 : _GEN_4873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4876 = ~io_inputBit ? 1'h0 : _GEN_4875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4877 = i == 10'h14 ? _GEN_4876 : _GEN_4875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4878 = io_inputBit ? 1'h0 : _GEN_4877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4879 = i == 10'h17 ? _GEN_4878 : _GEN_4877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4880 = ~io_inputBit ? 1'h0 : _GEN_4879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4881 = i == 10'h55 ? _GEN_4880 : _GEN_4879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4882 = ~io_inputBit | _GEN_4881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4883 = i == 10'h56 ? _GEN_4882 : _GEN_4881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4884 = ~io_inputBit ? 1'h0 : _GEN_4883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4885 = i == 10'h57 ? _GEN_4884 : _GEN_4883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4886 = ~io_inputBit | _GEN_4885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4887 = i == 10'h58 ? _GEN_4886 : _GEN_4885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4888 = ~io_inputBit ? 1'h0 : _GEN_4887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4889 = i == 10'h59 ? _GEN_4888 : _GEN_4887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4890 = ~io_inputBit | _GEN_4889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4891 = i == 10'h5a ? _GEN_4890 : _GEN_4889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4892 = io_inputBit | _GEN_4891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4893 = i == 10'h5b ? _GEN_4892 : _GEN_4891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4894 = io_inputBit ? 1'h0 : _GEN_4893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4895 = i == 10'h5c ? _GEN_4894 : _GEN_4893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4896 = io_inputBit | _GEN_4895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4897 = i == 10'h5d ? _GEN_4896 : _GEN_4895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4898 = io_inputBit ? 1'h0 : _GEN_4897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4899 = i == 10'h5e ? _GEN_4898 : _GEN_4897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4900 = io_inputBit | _GEN_4899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4901 = i == 10'h5f ? _GEN_4900 : _GEN_4899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4902 = io_inputBit ? 1'h0 : _GEN_4901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4903 = i == 10'h60 ? _GEN_4902 : _GEN_4901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4904 = ~io_inputBit ? 1'h0 : _GEN_4903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4905 = i == 10'hac ? _GEN_4904 : _GEN_4903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4906 = ~io_inputBit | _GEN_4905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4907 = i == 10'hae ? _GEN_4906 : _GEN_4905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4908 = ~io_inputBit ? 1'h0 : _GEN_4907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4909 = i == 10'hb0 ? _GEN_4908 : _GEN_4907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4910 = ~io_inputBit | _GEN_4909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4911 = i == 10'hb2 ? _GEN_4910 : _GEN_4909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4912 = ~io_inputBit ? 1'h0 : _GEN_4911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4913 = i == 10'hb4 ? _GEN_4912 : _GEN_4911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4914 = ~io_inputBit | _GEN_4913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4915 = i == 10'hb6 ? _GEN_4914 : _GEN_4913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4916 = ~io_inputBit ? 1'h0 : _GEN_4915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4917 = i == 10'hb7 ? _GEN_4916 : _GEN_4915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4918 = ~io_inputBit | _GEN_4917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4919 = i == 10'hb9 ? _GEN_4918 : _GEN_4917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4920 = ~io_inputBit ? 1'h0 : _GEN_4919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4921 = i == 10'hbb ? _GEN_4920 : _GEN_4919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4922 = ~io_inputBit | _GEN_4921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4923 = i == 10'hbd ? _GEN_4922 : _GEN_4921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4924 = ~io_inputBit ? 1'h0 : _GEN_4923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4925 = i == 10'hbf ? _GEN_4924 : _GEN_4923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4926 = ~io_inputBit | _GEN_4925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4927 = i == 10'hc1 ? _GEN_4926 : _GEN_4925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4928 = ~io_inputBit ? 1'h0 : _GEN_4927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4929 = i == 10'h15a ? _GEN_4928 : _GEN_4927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4930 = io_inputBit | _GEN_4929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4931 = i == 10'h15a ? _GEN_4930 : _GEN_4929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4932 = ~io_inputBit | _GEN_4931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4933 = i == 10'h15e ? _GEN_4932 : _GEN_4931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4934 = io_inputBit ? 1'h0 : _GEN_4933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4935 = i == 10'h15e ? _GEN_4934 : _GEN_4933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4936 = ~io_inputBit ? 1'h0 : _GEN_4935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4937 = i == 10'h162 ? _GEN_4936 : _GEN_4935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4938 = io_inputBit | _GEN_4937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4939 = i == 10'h162 ? _GEN_4938 : _GEN_4937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4940 = ~io_inputBit | _GEN_4939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4941 = i == 10'h166 ? _GEN_4940 : _GEN_4939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4942 = io_inputBit ? 1'h0 : _GEN_4941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4943 = i == 10'h166 ? _GEN_4942 : _GEN_4941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4944 = ~io_inputBit ? 1'h0 : _GEN_4943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4945 = i == 10'h16a ? _GEN_4944 : _GEN_4943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4946 = io_inputBit | _GEN_4945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4947 = i == 10'h16a ? _GEN_4946 : _GEN_4945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4948 = ~io_inputBit | _GEN_4947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4949 = i == 10'h16e ? _GEN_4948 : _GEN_4947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4950 = io_inputBit ? 1'h0 : _GEN_4949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4951 = i == 10'h16e ? _GEN_4950 : _GEN_4949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4952 = ~io_inputBit ? 1'h0 : _GEN_4951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4953 = i == 10'h170 ? _GEN_4952 : _GEN_4951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4954 = ~io_inputBit | _GEN_4953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4955 = i == 10'h174 ? _GEN_4954 : _GEN_4953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4956 = ~io_inputBit ? 1'h0 : _GEN_4955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4957 = i == 10'h178 ? _GEN_4956 : _GEN_4955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4958 = ~io_inputBit | _GEN_4957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4959 = i == 10'h17c ? _GEN_4958 : _GEN_4957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4960 = ~io_inputBit ? 1'h0 : _GEN_4959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4961 = i == 10'h180 ? _GEN_4960 : _GEN_4959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4962 = ~io_inputBit | _GEN_4961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4963 = i == 10'h184 ? _GEN_4962 : _GEN_4961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4964 = ~io_inputBit ? 1'h0 : _GEN_4963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4965 = i == 10'h2e2 ? _GEN_4964 : _GEN_4963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4966 = io_inputBit | _GEN_4965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4967 = i == 10'h2e2 ? _GEN_4966 : _GEN_4965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4968 = ~io_inputBit | _GEN_4967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4969 = i == 10'h2ea ? _GEN_4968 : _GEN_4967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4970 = io_inputBit ? 1'h0 : _GEN_4969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4971 = i == 10'h2ea ? _GEN_4970 : _GEN_4969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4972 = ~io_inputBit ? 1'h0 : _GEN_4971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4973 = i == 10'h2f2 ? _GEN_4972 : _GEN_4971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4974 = io_inputBit | _GEN_4973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4975 = i == 10'h2f2 ? _GEN_4974 : _GEN_4973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4976 = ~io_inputBit | _GEN_4975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4977 = i == 10'h2fa ? _GEN_4976 : _GEN_4975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4978 = io_inputBit ? 1'h0 : _GEN_4977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4979 = i == 10'h2fa ? _GEN_4978 : _GEN_4977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4980 = ~io_inputBit ? 1'h0 : _GEN_4979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4981 = i == 10'h302 ? _GEN_4980 : _GEN_4979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4982 = io_inputBit | _GEN_4981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4983 = i == 10'h302 ? _GEN_4982 : _GEN_4981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4984 = ~io_inputBit | _GEN_4983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4985 = i == 10'h30a ? _GEN_4984 : _GEN_4983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4986 = io_inputBit ? 1'h0 : _GEN_4985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4987 = i == 10'h30a ? _GEN_4986 : _GEN_4985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4988 = ~io_inputBit ? 1'h0 : _GEN_4351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4989 = i == 10'h1 ? _GEN_4988 : _GEN_4351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4990 = io_inputBit ? 1'h0 : _GEN_4989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4991 = i == 10'h2 ? _GEN_4990 : _GEN_4989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4992 = io_inputBit ? 1'h0 : _GEN_4991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4993 = i == 10'h5 ? _GEN_4992 : _GEN_4991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4994 = ~io_inputBit ? 1'h0 : _GEN_4993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4995 = i == 10'h9 ? _GEN_4994 : _GEN_4993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4996 = io_inputBit ? 1'h0 : _GEN_4995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4997 = i == 10'hb ? _GEN_4996 : _GEN_4995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4998 = ~io_inputBit ? 1'h0 : _GEN_4997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_4999 = i == 10'h14 ? _GEN_4998 : _GEN_4997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5000 = io_inputBit ? 1'h0 : _GEN_4999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5001 = i == 10'h17 ? _GEN_5000 : _GEN_4999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5002 = ~io_inputBit ? 1'h0 : _GEN_5001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5003 = i == 10'hab ? _GEN_5002 : _GEN_5001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5004 = ~io_inputBit | _GEN_5003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5005 = i == 10'hac ? _GEN_5004 : _GEN_5003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5006 = ~io_inputBit ? 1'h0 : _GEN_5005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5007 = i == 10'had ? _GEN_5006 : _GEN_5005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5008 = ~io_inputBit | _GEN_5007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5009 = i == 10'hae ? _GEN_5008 : _GEN_5007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5010 = ~io_inputBit ? 1'h0 : _GEN_5009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5011 = i == 10'haf ? _GEN_5010 : _GEN_5009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5012 = ~io_inputBit | _GEN_5011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5013 = i == 10'hb0 ? _GEN_5012 : _GEN_5011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5014 = ~io_inputBit ? 1'h0 : _GEN_5013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5015 = i == 10'hb1 ? _GEN_5014 : _GEN_5013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5016 = ~io_inputBit | _GEN_5015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5017 = i == 10'hb2 ? _GEN_5016 : _GEN_5015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5018 = ~io_inputBit ? 1'h0 : _GEN_5017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5019 = i == 10'hb3 ? _GEN_5018 : _GEN_5017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5020 = ~io_inputBit | _GEN_5019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5021 = i == 10'hb4 ? _GEN_5020 : _GEN_5019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5022 = ~io_inputBit ? 1'h0 : _GEN_5021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5023 = i == 10'hb5 ? _GEN_5022 : _GEN_5021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5024 = ~io_inputBit | _GEN_5023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5025 = i == 10'hb6 ? _GEN_5024 : _GEN_5023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5026 = ~io_inputBit ? 1'h0 : _GEN_5025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5027 = i == 10'hb7 ? _GEN_5026 : _GEN_5025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5028 = ~io_inputBit | _GEN_5027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5029 = i == 10'hb8 ? _GEN_5028 : _GEN_5027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5030 = ~io_inputBit ? 1'h0 : _GEN_5029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5031 = i == 10'hb9 ? _GEN_5030 : _GEN_5029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5032 = ~io_inputBit | _GEN_5031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5033 = i == 10'hba ? _GEN_5032 : _GEN_5031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5034 = ~io_inputBit ? 1'h0 : _GEN_5033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5035 = i == 10'hbb ? _GEN_5034 : _GEN_5033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5036 = ~io_inputBit | _GEN_5035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5037 = i == 10'hbc ? _GEN_5036 : _GEN_5035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5038 = ~io_inputBit ? 1'h0 : _GEN_5037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5039 = i == 10'hbd ? _GEN_5038 : _GEN_5037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5040 = ~io_inputBit | _GEN_5039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5041 = i == 10'hbe ? _GEN_5040 : _GEN_5039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5042 = ~io_inputBit ? 1'h0 : _GEN_5041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5043 = i == 10'hbf ? _GEN_5042 : _GEN_5041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5044 = ~io_inputBit | _GEN_5043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5045 = i == 10'hc0 ? _GEN_5044 : _GEN_5043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5046 = ~io_inputBit ? 1'h0 : _GEN_5045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5047 = i == 10'hc1 ? _GEN_5046 : _GEN_5045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5048 = ~io_inputBit | _GEN_5047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5049 = i == 10'hc2 ? _GEN_5048 : _GEN_5047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5050 = ~io_inputBit ? 1'h0 : _GEN_5049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5051 = i == 10'h158 ? _GEN_5050 : _GEN_5049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5052 = io_inputBit | _GEN_5051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5053 = i == 10'h158 ? _GEN_5052 : _GEN_5051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5054 = ~io_inputBit | _GEN_5053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5055 = i == 10'h15a ? _GEN_5054 : _GEN_5053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5056 = io_inputBit ? 1'h0 : _GEN_5055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5057 = i == 10'h15a ? _GEN_5056 : _GEN_5055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5058 = ~io_inputBit ? 1'h0 : _GEN_5057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5059 = i == 10'h15c ? _GEN_5058 : _GEN_5057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5060 = io_inputBit | _GEN_5059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5061 = i == 10'h15c ? _GEN_5060 : _GEN_5059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5062 = ~io_inputBit | _GEN_5061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5063 = i == 10'h15e ? _GEN_5062 : _GEN_5061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5064 = io_inputBit ? 1'h0 : _GEN_5063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5065 = i == 10'h15e ? _GEN_5064 : _GEN_5063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5066 = ~io_inputBit ? 1'h0 : _GEN_5065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5067 = i == 10'h160 ? _GEN_5066 : _GEN_5065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5068 = io_inputBit | _GEN_5067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5069 = i == 10'h160 ? _GEN_5068 : _GEN_5067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5070 = ~io_inputBit | _GEN_5069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5071 = i == 10'h162 ? _GEN_5070 : _GEN_5069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5072 = io_inputBit ? 1'h0 : _GEN_5071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5073 = i == 10'h162 ? _GEN_5072 : _GEN_5071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5074 = ~io_inputBit ? 1'h0 : _GEN_5073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5075 = i == 10'h164 ? _GEN_5074 : _GEN_5073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5076 = io_inputBit | _GEN_5075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5077 = i == 10'h164 ? _GEN_5076 : _GEN_5075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5078 = ~io_inputBit | _GEN_5077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5079 = i == 10'h166 ? _GEN_5078 : _GEN_5077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5080 = io_inputBit ? 1'h0 : _GEN_5079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5081 = i == 10'h166 ? _GEN_5080 : _GEN_5079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5082 = ~io_inputBit ? 1'h0 : _GEN_5081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5083 = i == 10'h168 ? _GEN_5082 : _GEN_5081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5084 = io_inputBit | _GEN_5083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5085 = i == 10'h168 ? _GEN_5084 : _GEN_5083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5086 = ~io_inputBit | _GEN_5085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5087 = i == 10'h16a ? _GEN_5086 : _GEN_5085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5088 = io_inputBit ? 1'h0 : _GEN_5087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5089 = i == 10'h16a ? _GEN_5088 : _GEN_5087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5090 = ~io_inputBit ? 1'h0 : _GEN_5089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5091 = i == 10'h16c ? _GEN_5090 : _GEN_5089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5092 = io_inputBit | _GEN_5091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5093 = i == 10'h16c ? _GEN_5092 : _GEN_5091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5094 = ~io_inputBit | _GEN_5093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5095 = i == 10'h16e ? _GEN_5094 : _GEN_5093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5096 = io_inputBit ? 1'h0 : _GEN_5095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5097 = i == 10'h16e ? _GEN_5096 : _GEN_5095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5098 = ~io_inputBit ? 1'h0 : _GEN_5097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5099 = i == 10'h170 ? _GEN_5098 : _GEN_5097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5100 = ~io_inputBit | _GEN_5099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5101 = i == 10'h172 ? _GEN_5100 : _GEN_5099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5102 = ~io_inputBit ? 1'h0 : _GEN_5101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5103 = i == 10'h174 ? _GEN_5102 : _GEN_5101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5104 = ~io_inputBit | _GEN_5103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5105 = i == 10'h176 ? _GEN_5104 : _GEN_5103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5106 = ~io_inputBit ? 1'h0 : _GEN_5105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5107 = i == 10'h178 ? _GEN_5106 : _GEN_5105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5108 = ~io_inputBit | _GEN_5107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5109 = i == 10'h17a ? _GEN_5108 : _GEN_5107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5110 = ~io_inputBit ? 1'h0 : _GEN_5109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5111 = i == 10'h17c ? _GEN_5110 : _GEN_5109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5112 = ~io_inputBit | _GEN_5111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5113 = i == 10'h17e ? _GEN_5112 : _GEN_5111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5114 = ~io_inputBit ? 1'h0 : _GEN_5113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5115 = i == 10'h180 ? _GEN_5114 : _GEN_5113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5116 = ~io_inputBit | _GEN_5115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5117 = i == 10'h182 ? _GEN_5116 : _GEN_5115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5118 = ~io_inputBit ? 1'h0 : _GEN_5117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5119 = i == 10'h184 ? _GEN_5118 : _GEN_5117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5120 = ~io_inputBit | _GEN_5119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5121 = i == 10'h186 ? _GEN_5120 : _GEN_5119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5122 = ~io_inputBit ? 1'h0 : _GEN_5121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5123 = i == 10'h2e2 ? _GEN_5122 : _GEN_5121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5124 = io_inputBit | _GEN_5123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5125 = i == 10'h2e2 ? _GEN_5124 : _GEN_5123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5126 = ~io_inputBit | _GEN_5125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5127 = i == 10'h2e6 ? _GEN_5126 : _GEN_5125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5128 = io_inputBit ? 1'h0 : _GEN_5127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5129 = i == 10'h2e6 ? _GEN_5128 : _GEN_5127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5130 = ~io_inputBit ? 1'h0 : _GEN_5129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5131 = i == 10'h2ea ? _GEN_5130 : _GEN_5129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5132 = io_inputBit | _GEN_5131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5133 = i == 10'h2ea ? _GEN_5132 : _GEN_5131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5134 = ~io_inputBit | _GEN_5133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5135 = i == 10'h2ee ? _GEN_5134 : _GEN_5133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5136 = io_inputBit ? 1'h0 : _GEN_5135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5137 = i == 10'h2ee ? _GEN_5136 : _GEN_5135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5138 = ~io_inputBit ? 1'h0 : _GEN_5137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5139 = i == 10'h2f2 ? _GEN_5138 : _GEN_5137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5140 = io_inputBit | _GEN_5139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5141 = i == 10'h2f2 ? _GEN_5140 : _GEN_5139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5142 = ~io_inputBit | _GEN_5141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5143 = i == 10'h2f6 ? _GEN_5142 : _GEN_5141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5144 = io_inputBit ? 1'h0 : _GEN_5143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5145 = i == 10'h2f6 ? _GEN_5144 : _GEN_5143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5146 = ~io_inputBit ? 1'h0 : _GEN_5145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5147 = i == 10'h2fa ? _GEN_5146 : _GEN_5145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5148 = io_inputBit | _GEN_5147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5149 = i == 10'h2fa ? _GEN_5148 : _GEN_5147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5150 = ~io_inputBit | _GEN_5149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5151 = i == 10'h2fe ? _GEN_5150 : _GEN_5149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5152 = io_inputBit ? 1'h0 : _GEN_5151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5153 = i == 10'h2fe ? _GEN_5152 : _GEN_5151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5154 = ~io_inputBit ? 1'h0 : _GEN_5153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5155 = i == 10'h302 ? _GEN_5154 : _GEN_5153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5156 = io_inputBit | _GEN_5155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5157 = i == 10'h302 ? _GEN_5156 : _GEN_5155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5158 = ~io_inputBit | _GEN_5157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5159 = i == 10'h306 ? _GEN_5158 : _GEN_5157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5160 = io_inputBit ? 1'h0 : _GEN_5159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5161 = i == 10'h306 ? _GEN_5160 : _GEN_5159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5162 = ~io_inputBit ? 1'h0 : _GEN_5161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5163 = i == 10'h30a ? _GEN_5162 : _GEN_5161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5164 = io_inputBit | _GEN_5163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5165 = i == 10'h30a ? _GEN_5164 : _GEN_5163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5166 = ~io_inputBit | _GEN_5165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5167 = i == 10'h30e ? _GEN_5166 : _GEN_5165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5168 = io_inputBit ? 1'h0 : _GEN_5167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5169 = i == 10'h30e ? _GEN_5168 : _GEN_5167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5170 = ~io_inputBit ? 1'h0 : _GEN_4421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5171 = i == 10'h1 ? _GEN_5170 : _GEN_4421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5172 = io_inputBit ? 1'h0 : _GEN_5171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5173 = i == 10'h2 ? _GEN_5172 : _GEN_5171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5174 = io_inputBit ? 1'h0 : _GEN_5173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5175 = i == 10'h5 ? _GEN_5174 : _GEN_5173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5176 = ~io_inputBit ? 1'h0 : _GEN_5175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5177 = i == 10'h9 ? _GEN_5176 : _GEN_5175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5178 = io_inputBit ? 1'h0 : _GEN_5177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5179 = i == 10'hb ? _GEN_5178 : _GEN_5177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5180 = ~io_inputBit ? 1'h0 : _GEN_5179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5181 = i == 10'h14 ? _GEN_5180 : _GEN_5179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5182 = io_inputBit ? 1'h0 : _GEN_5181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5183 = i == 10'h30 ? _GEN_5182 : _GEN_5181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5184 = io_inputBit ? 1'h0 : _GEN_5183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5185 = i == 10'h61 ? _GEN_5184 : _GEN_5183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5186 = io_inputBit ? 1'h0 : _GEN_5185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5187 = i == 10'hc3 ? _GEN_5186 : _GEN_5185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5188 = ~io_inputBit ? 1'h0 : _GEN_5187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5189 = i == 10'h157 ? _GEN_5188 : _GEN_5187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5190 = io_inputBit | _GEN_5189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5191 = i == 10'h157 ? _GEN_5190 : _GEN_5189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5192 = ~io_inputBit | _GEN_5191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5193 = i == 10'h158 ? _GEN_5192 : _GEN_5191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5194 = io_inputBit ? 1'h0 : _GEN_5193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5195 = i == 10'h158 ? _GEN_5194 : _GEN_5193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5196 = ~io_inputBit ? 1'h0 : _GEN_5195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5197 = i == 10'h159 ? _GEN_5196 : _GEN_5195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5198 = io_inputBit | _GEN_5197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5199 = i == 10'h159 ? _GEN_5198 : _GEN_5197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5200 = ~io_inputBit | _GEN_5199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5201 = i == 10'h15a ? _GEN_5200 : _GEN_5199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5202 = io_inputBit ? 1'h0 : _GEN_5201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5203 = i == 10'h15a ? _GEN_5202 : _GEN_5201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5204 = ~io_inputBit ? 1'h0 : _GEN_5203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5205 = i == 10'h15b ? _GEN_5204 : _GEN_5203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5206 = io_inputBit | _GEN_5205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5207 = i == 10'h15b ? _GEN_5206 : _GEN_5205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5208 = ~io_inputBit | _GEN_5207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5209 = i == 10'h15c ? _GEN_5208 : _GEN_5207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5210 = io_inputBit ? 1'h0 : _GEN_5209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5211 = i == 10'h15c ? _GEN_5210 : _GEN_5209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5212 = ~io_inputBit ? 1'h0 : _GEN_5211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5213 = i == 10'h15d ? _GEN_5212 : _GEN_5211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5214 = io_inputBit | _GEN_5213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5215 = i == 10'h15d ? _GEN_5214 : _GEN_5213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5216 = ~io_inputBit | _GEN_5215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5217 = i == 10'h15e ? _GEN_5216 : _GEN_5215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5218 = io_inputBit ? 1'h0 : _GEN_5217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5219 = i == 10'h15e ? _GEN_5218 : _GEN_5217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5220 = ~io_inputBit ? 1'h0 : _GEN_5219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5221 = i == 10'h15f ? _GEN_5220 : _GEN_5219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5222 = io_inputBit | _GEN_5221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5223 = i == 10'h15f ? _GEN_5222 : _GEN_5221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5224 = ~io_inputBit | _GEN_5223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5225 = i == 10'h160 ? _GEN_5224 : _GEN_5223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5226 = io_inputBit ? 1'h0 : _GEN_5225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5227 = i == 10'h160 ? _GEN_5226 : _GEN_5225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5228 = ~io_inputBit ? 1'h0 : _GEN_5227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5229 = i == 10'h161 ? _GEN_5228 : _GEN_5227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5230 = io_inputBit | _GEN_5229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5231 = i == 10'h161 ? _GEN_5230 : _GEN_5229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5232 = ~io_inputBit | _GEN_5231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5233 = i == 10'h162 ? _GEN_5232 : _GEN_5231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5234 = io_inputBit ? 1'h0 : _GEN_5233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5235 = i == 10'h162 ? _GEN_5234 : _GEN_5233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5236 = ~io_inputBit ? 1'h0 : _GEN_5235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5237 = i == 10'h163 ? _GEN_5236 : _GEN_5235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5238 = io_inputBit | _GEN_5237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5239 = i == 10'h163 ? _GEN_5238 : _GEN_5237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5240 = ~io_inputBit | _GEN_5239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5241 = i == 10'h164 ? _GEN_5240 : _GEN_5239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5242 = io_inputBit ? 1'h0 : _GEN_5241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5243 = i == 10'h164 ? _GEN_5242 : _GEN_5241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5244 = ~io_inputBit ? 1'h0 : _GEN_5243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5245 = i == 10'h165 ? _GEN_5244 : _GEN_5243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5246 = io_inputBit | _GEN_5245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5247 = i == 10'h165 ? _GEN_5246 : _GEN_5245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5248 = ~io_inputBit | _GEN_5247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5249 = i == 10'h166 ? _GEN_5248 : _GEN_5247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5250 = io_inputBit ? 1'h0 : _GEN_5249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5251 = i == 10'h166 ? _GEN_5250 : _GEN_5249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5252 = ~io_inputBit ? 1'h0 : _GEN_5251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5253 = i == 10'h167 ? _GEN_5252 : _GEN_5251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5254 = io_inputBit | _GEN_5253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5255 = i == 10'h167 ? _GEN_5254 : _GEN_5253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5256 = ~io_inputBit | _GEN_5255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5257 = i == 10'h168 ? _GEN_5256 : _GEN_5255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5258 = io_inputBit ? 1'h0 : _GEN_5257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5259 = i == 10'h168 ? _GEN_5258 : _GEN_5257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5260 = ~io_inputBit ? 1'h0 : _GEN_5259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5261 = i == 10'h169 ? _GEN_5260 : _GEN_5259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5262 = io_inputBit | _GEN_5261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5263 = i == 10'h169 ? _GEN_5262 : _GEN_5261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5264 = ~io_inputBit | _GEN_5263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5265 = i == 10'h16a ? _GEN_5264 : _GEN_5263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5266 = io_inputBit ? 1'h0 : _GEN_5265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5267 = i == 10'h16a ? _GEN_5266 : _GEN_5265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5268 = ~io_inputBit ? 1'h0 : _GEN_5267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5269 = i == 10'h16b ? _GEN_5268 : _GEN_5267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5270 = io_inputBit | _GEN_5269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5271 = i == 10'h16b ? _GEN_5270 : _GEN_5269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5272 = ~io_inputBit | _GEN_5271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5273 = i == 10'h16c ? _GEN_5272 : _GEN_5271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5274 = io_inputBit ? 1'h0 : _GEN_5273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5275 = i == 10'h16c ? _GEN_5274 : _GEN_5273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5276 = ~io_inputBit ? 1'h0 : _GEN_5275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5277 = i == 10'h16d ? _GEN_5276 : _GEN_5275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5278 = io_inputBit | _GEN_5277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5279 = i == 10'h16d ? _GEN_5278 : _GEN_5277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5280 = ~io_inputBit | _GEN_5279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5281 = i == 10'h16e ? _GEN_5280 : _GEN_5279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5282 = io_inputBit ? 1'h0 : _GEN_5281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5283 = i == 10'h16e ? _GEN_5282 : _GEN_5281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5284 = ~io_inputBit ? 1'h0 : _GEN_5283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5285 = i == 10'h16f ? _GEN_5284 : _GEN_5283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5286 = ~io_inputBit ? 1'h0 : _GEN_5285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5287 = i == 10'h170 ? _GEN_5286 : _GEN_5285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5288 = ~io_inputBit | _GEN_5287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5289 = i == 10'h171 ? _GEN_5288 : _GEN_5287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5290 = ~io_inputBit ? 1'h0 : _GEN_5289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5291 = i == 10'h172 ? _GEN_5290 : _GEN_5289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5292 = ~io_inputBit | _GEN_5291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5293 = i == 10'h173 ? _GEN_5292 : _GEN_5291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5294 = ~io_inputBit ? 1'h0 : _GEN_5293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5295 = i == 10'h174 ? _GEN_5294 : _GEN_5293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5296 = ~io_inputBit | _GEN_5295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5297 = i == 10'h175 ? _GEN_5296 : _GEN_5295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5298 = ~io_inputBit ? 1'h0 : _GEN_5297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5299 = i == 10'h176 ? _GEN_5298 : _GEN_5297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5300 = ~io_inputBit | _GEN_5299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5301 = i == 10'h177 ? _GEN_5300 : _GEN_5299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5302 = ~io_inputBit ? 1'h0 : _GEN_5301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5303 = i == 10'h178 ? _GEN_5302 : _GEN_5301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5304 = ~io_inputBit | _GEN_5303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5305 = i == 10'h179 ? _GEN_5304 : _GEN_5303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5306 = ~io_inputBit ? 1'h0 : _GEN_5305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5307 = i == 10'h17a ? _GEN_5306 : _GEN_5305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5308 = ~io_inputBit | _GEN_5307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5309 = i == 10'h17b ? _GEN_5308 : _GEN_5307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5310 = ~io_inputBit ? 1'h0 : _GEN_5309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5311 = i == 10'h17c ? _GEN_5310 : _GEN_5309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5312 = ~io_inputBit | _GEN_5311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5313 = i == 10'h17d ? _GEN_5312 : _GEN_5311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5314 = ~io_inputBit ? 1'h0 : _GEN_5313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5315 = i == 10'h17e ? _GEN_5314 : _GEN_5313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5316 = ~io_inputBit | _GEN_5315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5317 = i == 10'h17f ? _GEN_5316 : _GEN_5315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5318 = ~io_inputBit ? 1'h0 : _GEN_5317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5319 = i == 10'h180 ? _GEN_5318 : _GEN_5317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5320 = ~io_inputBit | _GEN_5319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5321 = i == 10'h181 ? _GEN_5320 : _GEN_5319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5322 = ~io_inputBit ? 1'h0 : _GEN_5321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5323 = i == 10'h182 ? _GEN_5322 : _GEN_5321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5324 = ~io_inputBit | _GEN_5323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5325 = i == 10'h183 ? _GEN_5324 : _GEN_5323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5326 = ~io_inputBit ? 1'h0 : _GEN_5325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5327 = i == 10'h184 ? _GEN_5326 : _GEN_5325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5328 = ~io_inputBit | _GEN_5327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5329 = i == 10'h185 ? _GEN_5328 : _GEN_5327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5330 = ~io_inputBit ? 1'h0 : _GEN_5329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5331 = i == 10'h186 ? _GEN_5330 : _GEN_5329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5332 = ~io_inputBit | _GEN_5331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5333 = i == 10'h187 ? _GEN_5332 : _GEN_5331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5334 = ~io_inputBit | _GEN_5333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5335 = i == 10'h2e0 ? _GEN_5334 : _GEN_5333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5336 = io_inputBit ? 1'h0 : _GEN_5335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5337 = i == 10'h2e0 ? _GEN_5336 : _GEN_5335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5338 = ~io_inputBit ? 1'h0 : _GEN_5337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5339 = i == 10'h2e2 ? _GEN_5338 : _GEN_5337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5340 = io_inputBit | _GEN_5339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5341 = i == 10'h2e2 ? _GEN_5340 : _GEN_5339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5342 = ~io_inputBit | _GEN_5341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5343 = i == 10'h2e4 ? _GEN_5342 : _GEN_5341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5344 = io_inputBit ? 1'h0 : _GEN_5343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5345 = i == 10'h2e4 ? _GEN_5344 : _GEN_5343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5346 = ~io_inputBit ? 1'h0 : _GEN_5345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5347 = i == 10'h2e6 ? _GEN_5346 : _GEN_5345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5348 = io_inputBit | _GEN_5347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5349 = i == 10'h2e6 ? _GEN_5348 : _GEN_5347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5350 = ~io_inputBit | _GEN_5349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5351 = i == 10'h2e8 ? _GEN_5350 : _GEN_5349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5352 = io_inputBit ? 1'h0 : _GEN_5351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5353 = i == 10'h2e8 ? _GEN_5352 : _GEN_5351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5354 = ~io_inputBit ? 1'h0 : _GEN_5353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5355 = i == 10'h2ea ? _GEN_5354 : _GEN_5353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5356 = io_inputBit | _GEN_5355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5357 = i == 10'h2ea ? _GEN_5356 : _GEN_5355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5358 = ~io_inputBit | _GEN_5357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5359 = i == 10'h2ec ? _GEN_5358 : _GEN_5357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5360 = io_inputBit ? 1'h0 : _GEN_5359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5361 = i == 10'h2ec ? _GEN_5360 : _GEN_5359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5362 = ~io_inputBit ? 1'h0 : _GEN_5361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5363 = i == 10'h2ee ? _GEN_5362 : _GEN_5361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5364 = io_inputBit | _GEN_5363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5365 = i == 10'h2ee ? _GEN_5364 : _GEN_5363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5366 = ~io_inputBit | _GEN_5365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5367 = i == 10'h2f0 ? _GEN_5366 : _GEN_5365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5368 = io_inputBit ? 1'h0 : _GEN_5367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5369 = i == 10'h2f0 ? _GEN_5368 : _GEN_5367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5370 = ~io_inputBit ? 1'h0 : _GEN_5369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5371 = i == 10'h2f2 ? _GEN_5370 : _GEN_5369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5372 = io_inputBit | _GEN_5371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5373 = i == 10'h2f2 ? _GEN_5372 : _GEN_5371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5374 = ~io_inputBit | _GEN_5373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5375 = i == 10'h2f4 ? _GEN_5374 : _GEN_5373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5376 = io_inputBit ? 1'h0 : _GEN_5375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5377 = i == 10'h2f4 ? _GEN_5376 : _GEN_5375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5378 = ~io_inputBit ? 1'h0 : _GEN_5377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5379 = i == 10'h2f6 ? _GEN_5378 : _GEN_5377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5380 = io_inputBit | _GEN_5379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5381 = i == 10'h2f6 ? _GEN_5380 : _GEN_5379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5382 = ~io_inputBit | _GEN_5381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5383 = i == 10'h2f8 ? _GEN_5382 : _GEN_5381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5384 = io_inputBit ? 1'h0 : _GEN_5383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5385 = i == 10'h2f8 ? _GEN_5384 : _GEN_5383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5386 = ~io_inputBit ? 1'h0 : _GEN_5385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5387 = i == 10'h2fa ? _GEN_5386 : _GEN_5385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5388 = io_inputBit | _GEN_5387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5389 = i == 10'h2fa ? _GEN_5388 : _GEN_5387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5390 = ~io_inputBit | _GEN_5389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5391 = i == 10'h2fc ? _GEN_5390 : _GEN_5389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5392 = io_inputBit ? 1'h0 : _GEN_5391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5393 = i == 10'h2fc ? _GEN_5392 : _GEN_5391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5394 = ~io_inputBit ? 1'h0 : _GEN_5393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5395 = i == 10'h2fe ? _GEN_5394 : _GEN_5393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5396 = io_inputBit | _GEN_5395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5397 = i == 10'h2fe ? _GEN_5396 : _GEN_5395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5398 = ~io_inputBit | _GEN_5397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5399 = i == 10'h300 ? _GEN_5398 : _GEN_5397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5400 = io_inputBit ? 1'h0 : _GEN_5399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5401 = i == 10'h300 ? _GEN_5400 : _GEN_5399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5402 = ~io_inputBit ? 1'h0 : _GEN_5401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5403 = i == 10'h302 ? _GEN_5402 : _GEN_5401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5404 = io_inputBit | _GEN_5403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5405 = i == 10'h302 ? _GEN_5404 : _GEN_5403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5406 = ~io_inputBit | _GEN_5405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5407 = i == 10'h304 ? _GEN_5406 : _GEN_5405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5408 = io_inputBit ? 1'h0 : _GEN_5407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5409 = i == 10'h304 ? _GEN_5408 : _GEN_5407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5410 = ~io_inputBit ? 1'h0 : _GEN_5409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5411 = i == 10'h306 ? _GEN_5410 : _GEN_5409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5412 = io_inputBit | _GEN_5411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5413 = i == 10'h306 ? _GEN_5412 : _GEN_5411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5414 = ~io_inputBit | _GEN_5413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5415 = i == 10'h308 ? _GEN_5414 : _GEN_5413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5416 = io_inputBit ? 1'h0 : _GEN_5415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5417 = i == 10'h308 ? _GEN_5416 : _GEN_5415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5418 = ~io_inputBit ? 1'h0 : _GEN_5417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5419 = i == 10'h30a ? _GEN_5418 : _GEN_5417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5420 = io_inputBit | _GEN_5419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5421 = i == 10'h30a ? _GEN_5420 : _GEN_5419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5422 = ~io_inputBit | _GEN_5421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5423 = i == 10'h30c ? _GEN_5422 : _GEN_5421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5424 = io_inputBit ? 1'h0 : _GEN_5423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5425 = i == 10'h30c ? _GEN_5424 : _GEN_5423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5426 = ~io_inputBit ? 1'h0 : _GEN_5425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5427 = i == 10'h30e ? _GEN_5426 : _GEN_5425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5428 = io_inputBit | _GEN_5427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5429 = i == 10'h30e ? _GEN_5428 : _GEN_5427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5430 = ~io_inputBit | _GEN_5429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5431 = i == 10'h310 ? _GEN_5430 : _GEN_5429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5432 = io_inputBit ? 1'h0 : _GEN_5431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5433 = i == 10'h310 ? _GEN_5432 : _GEN_5431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5434 = ~io_inputBit ? 1'h0 : _GEN_4537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5435 = i == 10'h1 ? _GEN_5434 : _GEN_4537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5436 = io_inputBit ? 1'h0 : _GEN_5435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5437 = i == 10'h2 ? _GEN_5436 : _GEN_5435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5438 = io_inputBit ? 1'h0 : _GEN_5437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5439 = i == 10'h5 ? _GEN_5438 : _GEN_5437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5440 = ~io_inputBit ? 1'h0 : _GEN_5439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5441 = i == 10'h9 ? _GEN_5440 : _GEN_5439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5442 = io_inputBit ? 1'h0 : _GEN_5441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5443 = i == 10'hb ? _GEN_5442 : _GEN_5441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5444 = ~io_inputBit ? 1'h0 : _GEN_5443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5445 = i == 10'h14 ? _GEN_5444 : _GEN_5443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5446 = io_inputBit ? 1'h0 : _GEN_5445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5447 = i == 10'h30 ? _GEN_5446 : _GEN_5445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5448 = io_inputBit ? 1'h0 : _GEN_5447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5449 = i == 10'h61 ? _GEN_5448 : _GEN_5447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5450 = ~io_inputBit | _GEN_5449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5451 = i == 10'h157 ? _GEN_5450 : _GEN_5449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5452 = io_inputBit ? 1'h0 : _GEN_5451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5453 = i == 10'h157 ? _GEN_5452 : _GEN_5451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5454 = ~io_inputBit | _GEN_5453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5455 = i == 10'h158 ? _GEN_5454 : _GEN_5453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5456 = io_inputBit ? 1'h0 : _GEN_5455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5457 = i == 10'h158 ? _GEN_5456 : _GEN_5455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5458 = ~io_inputBit | _GEN_5457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5459 = i == 10'h159 ? _GEN_5458 : _GEN_5457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5460 = io_inputBit ? 1'h0 : _GEN_5459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5461 = i == 10'h159 ? _GEN_5460 : _GEN_5459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5462 = ~io_inputBit | _GEN_5461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5463 = i == 10'h15a ? _GEN_5462 : _GEN_5461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5464 = io_inputBit ? 1'h0 : _GEN_5463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5465 = i == 10'h15a ? _GEN_5464 : _GEN_5463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5466 = ~io_inputBit | _GEN_5465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5467 = i == 10'h15b ? _GEN_5466 : _GEN_5465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5468 = io_inputBit ? 1'h0 : _GEN_5467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5469 = i == 10'h15b ? _GEN_5468 : _GEN_5467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5470 = ~io_inputBit | _GEN_5469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5471 = i == 10'h15c ? _GEN_5470 : _GEN_5469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5472 = io_inputBit ? 1'h0 : _GEN_5471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5473 = i == 10'h15c ? _GEN_5472 : _GEN_5471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5474 = ~io_inputBit | _GEN_5473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5475 = i == 10'h15d ? _GEN_5474 : _GEN_5473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5476 = io_inputBit ? 1'h0 : _GEN_5475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5477 = i == 10'h15d ? _GEN_5476 : _GEN_5475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5478 = ~io_inputBit | _GEN_5477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5479 = i == 10'h15e ? _GEN_5478 : _GEN_5477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5480 = io_inputBit ? 1'h0 : _GEN_5479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5481 = i == 10'h15e ? _GEN_5480 : _GEN_5479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5482 = ~io_inputBit | _GEN_5481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5483 = i == 10'h15f ? _GEN_5482 : _GEN_5481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5484 = io_inputBit ? 1'h0 : _GEN_5483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5485 = i == 10'h15f ? _GEN_5484 : _GEN_5483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5486 = ~io_inputBit | _GEN_5485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5487 = i == 10'h160 ? _GEN_5486 : _GEN_5485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5488 = io_inputBit ? 1'h0 : _GEN_5487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5489 = i == 10'h160 ? _GEN_5488 : _GEN_5487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5490 = ~io_inputBit | _GEN_5489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5491 = i == 10'h161 ? _GEN_5490 : _GEN_5489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5492 = io_inputBit ? 1'h0 : _GEN_5491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5493 = i == 10'h161 ? _GEN_5492 : _GEN_5491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5494 = ~io_inputBit | _GEN_5493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5495 = i == 10'h162 ? _GEN_5494 : _GEN_5493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5496 = io_inputBit ? 1'h0 : _GEN_5495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5497 = i == 10'h162 ? _GEN_5496 : _GEN_5495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5498 = ~io_inputBit | _GEN_5497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5499 = i == 10'h163 ? _GEN_5498 : _GEN_5497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5500 = io_inputBit ? 1'h0 : _GEN_5499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5501 = i == 10'h163 ? _GEN_5500 : _GEN_5499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5502 = ~io_inputBit | _GEN_5501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5503 = i == 10'h164 ? _GEN_5502 : _GEN_5501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5504 = io_inputBit ? 1'h0 : _GEN_5503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5505 = i == 10'h164 ? _GEN_5504 : _GEN_5503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5506 = ~io_inputBit | _GEN_5505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5507 = i == 10'h165 ? _GEN_5506 : _GEN_5505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5508 = io_inputBit ? 1'h0 : _GEN_5507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5509 = i == 10'h165 ? _GEN_5508 : _GEN_5507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5510 = ~io_inputBit | _GEN_5509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5511 = i == 10'h166 ? _GEN_5510 : _GEN_5509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5512 = io_inputBit ? 1'h0 : _GEN_5511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5513 = i == 10'h166 ? _GEN_5512 : _GEN_5511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5514 = ~io_inputBit | _GEN_5513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5515 = i == 10'h167 ? _GEN_5514 : _GEN_5513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5516 = io_inputBit ? 1'h0 : _GEN_5515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5517 = i == 10'h167 ? _GEN_5516 : _GEN_5515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5518 = ~io_inputBit | _GEN_5517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5519 = i == 10'h168 ? _GEN_5518 : _GEN_5517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5520 = io_inputBit ? 1'h0 : _GEN_5519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5521 = i == 10'h168 ? _GEN_5520 : _GEN_5519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5522 = ~io_inputBit | _GEN_5521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5523 = i == 10'h169 ? _GEN_5522 : _GEN_5521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5524 = io_inputBit ? 1'h0 : _GEN_5523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5525 = i == 10'h169 ? _GEN_5524 : _GEN_5523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5526 = ~io_inputBit | _GEN_5525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5527 = i == 10'h16a ? _GEN_5526 : _GEN_5525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5528 = io_inputBit ? 1'h0 : _GEN_5527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5529 = i == 10'h16a ? _GEN_5528 : _GEN_5527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5530 = ~io_inputBit | _GEN_5529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5531 = i == 10'h16b ? _GEN_5530 : _GEN_5529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5532 = io_inputBit ? 1'h0 : _GEN_5531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5533 = i == 10'h16b ? _GEN_5532 : _GEN_5531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5534 = ~io_inputBit | _GEN_5533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5535 = i == 10'h16c ? _GEN_5534 : _GEN_5533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5536 = io_inputBit ? 1'h0 : _GEN_5535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5537 = i == 10'h16c ? _GEN_5536 : _GEN_5535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5538 = ~io_inputBit | _GEN_5537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5539 = i == 10'h16d ? _GEN_5538 : _GEN_5537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5540 = io_inputBit ? 1'h0 : _GEN_5539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5541 = i == 10'h16d ? _GEN_5540 : _GEN_5539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5542 = ~io_inputBit | _GEN_5541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5543 = i == 10'h16e ? _GEN_5542 : _GEN_5541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5544 = io_inputBit ? 1'h0 : _GEN_5543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5545 = i == 10'h16e ? _GEN_5544 : _GEN_5543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5546 = ~io_inputBit | _GEN_5545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5547 = i == 10'h16f ? _GEN_5546 : _GEN_5545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5548 = io_inputBit ? 1'h0 : _GEN_5547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5549 = i == 10'h188 ? _GEN_5548 : _GEN_5547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5550 = ~io_inputBit ? 1'h0 : _GEN_5549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5551 = i == 10'h2e0 ? _GEN_5550 : _GEN_5549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5552 = io_inputBit | _GEN_5551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5553 = i == 10'h2e0 ? _GEN_5552 : _GEN_5551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5554 = ~io_inputBit | _GEN_5553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5555 = i == 10'h2e1 ? _GEN_5554 : _GEN_5553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5556 = io_inputBit ? 1'h0 : _GEN_5555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5557 = i == 10'h2e1 ? _GEN_5556 : _GEN_5555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5558 = ~io_inputBit ? 1'h0 : _GEN_5557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5559 = i == 10'h2e2 ? _GEN_5558 : _GEN_5557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5560 = io_inputBit | _GEN_5559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5561 = i == 10'h2e2 ? _GEN_5560 : _GEN_5559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5562 = ~io_inputBit | _GEN_5561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5563 = i == 10'h2e3 ? _GEN_5562 : _GEN_5561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5564 = io_inputBit ? 1'h0 : _GEN_5563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5565 = i == 10'h2e3 ? _GEN_5564 : _GEN_5563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5566 = ~io_inputBit ? 1'h0 : _GEN_5565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5567 = i == 10'h2e4 ? _GEN_5566 : _GEN_5565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5568 = io_inputBit | _GEN_5567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5569 = i == 10'h2e4 ? _GEN_5568 : _GEN_5567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5570 = ~io_inputBit | _GEN_5569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5571 = i == 10'h2e5 ? _GEN_5570 : _GEN_5569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5572 = io_inputBit ? 1'h0 : _GEN_5571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5573 = i == 10'h2e5 ? _GEN_5572 : _GEN_5571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5574 = ~io_inputBit ? 1'h0 : _GEN_5573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5575 = i == 10'h2e6 ? _GEN_5574 : _GEN_5573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5576 = io_inputBit | _GEN_5575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5577 = i == 10'h2e6 ? _GEN_5576 : _GEN_5575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5578 = ~io_inputBit | _GEN_5577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5579 = i == 10'h2e7 ? _GEN_5578 : _GEN_5577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5580 = io_inputBit ? 1'h0 : _GEN_5579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5581 = i == 10'h2e7 ? _GEN_5580 : _GEN_5579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5582 = ~io_inputBit ? 1'h0 : _GEN_5581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5583 = i == 10'h2e8 ? _GEN_5582 : _GEN_5581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5584 = io_inputBit | _GEN_5583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5585 = i == 10'h2e8 ? _GEN_5584 : _GEN_5583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5586 = ~io_inputBit | _GEN_5585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5587 = i == 10'h2e9 ? _GEN_5586 : _GEN_5585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5588 = io_inputBit ? 1'h0 : _GEN_5587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5589 = i == 10'h2e9 ? _GEN_5588 : _GEN_5587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5590 = ~io_inputBit ? 1'h0 : _GEN_5589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5591 = i == 10'h2ea ? _GEN_5590 : _GEN_5589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5592 = io_inputBit | _GEN_5591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5593 = i == 10'h2ea ? _GEN_5592 : _GEN_5591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5594 = ~io_inputBit | _GEN_5593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5595 = i == 10'h2eb ? _GEN_5594 : _GEN_5593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5596 = io_inputBit ? 1'h0 : _GEN_5595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5597 = i == 10'h2eb ? _GEN_5596 : _GEN_5595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5598 = ~io_inputBit ? 1'h0 : _GEN_5597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5599 = i == 10'h2ec ? _GEN_5598 : _GEN_5597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5600 = io_inputBit | _GEN_5599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5601 = i == 10'h2ec ? _GEN_5600 : _GEN_5599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5602 = ~io_inputBit | _GEN_5601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5603 = i == 10'h2ed ? _GEN_5602 : _GEN_5601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5604 = io_inputBit ? 1'h0 : _GEN_5603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5605 = i == 10'h2ed ? _GEN_5604 : _GEN_5603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5606 = ~io_inputBit ? 1'h0 : _GEN_5605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5607 = i == 10'h2ee ? _GEN_5606 : _GEN_5605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5608 = io_inputBit | _GEN_5607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5609 = i == 10'h2ee ? _GEN_5608 : _GEN_5607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5610 = ~io_inputBit | _GEN_5609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5611 = i == 10'h2ef ? _GEN_5610 : _GEN_5609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5612 = io_inputBit ? 1'h0 : _GEN_5611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5613 = i == 10'h2ef ? _GEN_5612 : _GEN_5611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5614 = ~io_inputBit ? 1'h0 : _GEN_5613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5615 = i == 10'h2f0 ? _GEN_5614 : _GEN_5613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5616 = io_inputBit | _GEN_5615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5617 = i == 10'h2f0 ? _GEN_5616 : _GEN_5615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5618 = ~io_inputBit | _GEN_5617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5619 = i == 10'h2f1 ? _GEN_5618 : _GEN_5617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5620 = io_inputBit ? 1'h0 : _GEN_5619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5621 = i == 10'h2f1 ? _GEN_5620 : _GEN_5619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5622 = ~io_inputBit ? 1'h0 : _GEN_5621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5623 = i == 10'h2f2 ? _GEN_5622 : _GEN_5621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5624 = io_inputBit | _GEN_5623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5625 = i == 10'h2f2 ? _GEN_5624 : _GEN_5623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5626 = ~io_inputBit | _GEN_5625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5627 = i == 10'h2f3 ? _GEN_5626 : _GEN_5625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5628 = io_inputBit ? 1'h0 : _GEN_5627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5629 = i == 10'h2f3 ? _GEN_5628 : _GEN_5627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5630 = ~io_inputBit ? 1'h0 : _GEN_5629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5631 = i == 10'h2f4 ? _GEN_5630 : _GEN_5629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5632 = io_inputBit | _GEN_5631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5633 = i == 10'h2f4 ? _GEN_5632 : _GEN_5631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5634 = ~io_inputBit | _GEN_5633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5635 = i == 10'h2f5 ? _GEN_5634 : _GEN_5633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5636 = io_inputBit ? 1'h0 : _GEN_5635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5637 = i == 10'h2f5 ? _GEN_5636 : _GEN_5635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5638 = ~io_inputBit ? 1'h0 : _GEN_5637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5639 = i == 10'h2f6 ? _GEN_5638 : _GEN_5637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5640 = io_inputBit | _GEN_5639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5641 = i == 10'h2f6 ? _GEN_5640 : _GEN_5639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5642 = ~io_inputBit | _GEN_5641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5643 = i == 10'h2f7 ? _GEN_5642 : _GEN_5641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5644 = io_inputBit ? 1'h0 : _GEN_5643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5645 = i == 10'h2f7 ? _GEN_5644 : _GEN_5643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5646 = ~io_inputBit ? 1'h0 : _GEN_5645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5647 = i == 10'h2f8 ? _GEN_5646 : _GEN_5645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5648 = io_inputBit | _GEN_5647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5649 = i == 10'h2f8 ? _GEN_5648 : _GEN_5647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5650 = ~io_inputBit | _GEN_5649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5651 = i == 10'h2f9 ? _GEN_5650 : _GEN_5649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5652 = io_inputBit ? 1'h0 : _GEN_5651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5653 = i == 10'h2f9 ? _GEN_5652 : _GEN_5651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5654 = ~io_inputBit ? 1'h0 : _GEN_5653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5655 = i == 10'h2fa ? _GEN_5654 : _GEN_5653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5656 = io_inputBit | _GEN_5655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5657 = i == 10'h2fa ? _GEN_5656 : _GEN_5655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5658 = ~io_inputBit | _GEN_5657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5659 = i == 10'h2fb ? _GEN_5658 : _GEN_5657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5660 = io_inputBit ? 1'h0 : _GEN_5659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5661 = i == 10'h2fb ? _GEN_5660 : _GEN_5659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5662 = ~io_inputBit ? 1'h0 : _GEN_5661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5663 = i == 10'h2fc ? _GEN_5662 : _GEN_5661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5664 = io_inputBit | _GEN_5663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5665 = i == 10'h2fc ? _GEN_5664 : _GEN_5663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5666 = ~io_inputBit | _GEN_5665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5667 = i == 10'h2fd ? _GEN_5666 : _GEN_5665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5668 = io_inputBit ? 1'h0 : _GEN_5667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5669 = i == 10'h2fd ? _GEN_5668 : _GEN_5667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5670 = ~io_inputBit ? 1'h0 : _GEN_5669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5671 = i == 10'h2fe ? _GEN_5670 : _GEN_5669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5672 = io_inputBit | _GEN_5671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5673 = i == 10'h2fe ? _GEN_5672 : _GEN_5671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5674 = ~io_inputBit | _GEN_5673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5675 = i == 10'h2ff ? _GEN_5674 : _GEN_5673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5676 = io_inputBit ? 1'h0 : _GEN_5675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5677 = i == 10'h2ff ? _GEN_5676 : _GEN_5675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5678 = ~io_inputBit ? 1'h0 : _GEN_5677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5679 = i == 10'h300 ? _GEN_5678 : _GEN_5677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5680 = io_inputBit | _GEN_5679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5681 = i == 10'h300 ? _GEN_5680 : _GEN_5679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5682 = ~io_inputBit | _GEN_5681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5683 = i == 10'h301 ? _GEN_5682 : _GEN_5681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5684 = io_inputBit ? 1'h0 : _GEN_5683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5685 = i == 10'h301 ? _GEN_5684 : _GEN_5683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5686 = ~io_inputBit ? 1'h0 : _GEN_5685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5687 = i == 10'h302 ? _GEN_5686 : _GEN_5685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5688 = io_inputBit | _GEN_5687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5689 = i == 10'h302 ? _GEN_5688 : _GEN_5687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5690 = ~io_inputBit | _GEN_5689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5691 = i == 10'h303 ? _GEN_5690 : _GEN_5689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5692 = io_inputBit ? 1'h0 : _GEN_5691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5693 = i == 10'h303 ? _GEN_5692 : _GEN_5691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5694 = ~io_inputBit ? 1'h0 : _GEN_5693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5695 = i == 10'h304 ? _GEN_5694 : _GEN_5693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5696 = io_inputBit | _GEN_5695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5697 = i == 10'h304 ? _GEN_5696 : _GEN_5695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5698 = ~io_inputBit | _GEN_5697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5699 = i == 10'h305 ? _GEN_5698 : _GEN_5697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5700 = io_inputBit ? 1'h0 : _GEN_5699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5701 = i == 10'h305 ? _GEN_5700 : _GEN_5699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5702 = ~io_inputBit ? 1'h0 : _GEN_5701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5703 = i == 10'h306 ? _GEN_5702 : _GEN_5701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5704 = io_inputBit | _GEN_5703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5705 = i == 10'h306 ? _GEN_5704 : _GEN_5703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5706 = ~io_inputBit | _GEN_5705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5707 = i == 10'h307 ? _GEN_5706 : _GEN_5705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5708 = io_inputBit ? 1'h0 : _GEN_5707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5709 = i == 10'h307 ? _GEN_5708 : _GEN_5707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5710 = ~io_inputBit ? 1'h0 : _GEN_5709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5711 = i == 10'h308 ? _GEN_5710 : _GEN_5709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5712 = io_inputBit | _GEN_5711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5713 = i == 10'h308 ? _GEN_5712 : _GEN_5711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5714 = ~io_inputBit | _GEN_5713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5715 = i == 10'h309 ? _GEN_5714 : _GEN_5713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5716 = io_inputBit ? 1'h0 : _GEN_5715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5717 = i == 10'h309 ? _GEN_5716 : _GEN_5715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5718 = ~io_inputBit ? 1'h0 : _GEN_5717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5719 = i == 10'h30a ? _GEN_5718 : _GEN_5717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5720 = io_inputBit | _GEN_5719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5721 = i == 10'h30a ? _GEN_5720 : _GEN_5719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5722 = ~io_inputBit | _GEN_5721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5723 = i == 10'h30b ? _GEN_5722 : _GEN_5721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5724 = io_inputBit ? 1'h0 : _GEN_5723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5725 = i == 10'h30b ? _GEN_5724 : _GEN_5723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5726 = ~io_inputBit ? 1'h0 : _GEN_5725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5727 = i == 10'h30c ? _GEN_5726 : _GEN_5725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5728 = io_inputBit | _GEN_5727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5729 = i == 10'h30c ? _GEN_5728 : _GEN_5727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5730 = ~io_inputBit | _GEN_5729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5731 = i == 10'h30d ? _GEN_5730 : _GEN_5729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5732 = io_inputBit ? 1'h0 : _GEN_5731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5733 = i == 10'h30d ? _GEN_5732 : _GEN_5731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5734 = ~io_inputBit ? 1'h0 : _GEN_5733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5735 = i == 10'h30e ? _GEN_5734 : _GEN_5733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5736 = io_inputBit | _GEN_5735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5737 = i == 10'h30e ? _GEN_5736 : _GEN_5735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5738 = ~io_inputBit | _GEN_5737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5739 = i == 10'h30f ? _GEN_5738 : _GEN_5737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5740 = io_inputBit ? 1'h0 : _GEN_5739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5741 = i == 10'h30f ? _GEN_5740 : _GEN_5739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5742 = ~io_inputBit ? 1'h0 : _GEN_5741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5743 = i == 10'h310 ? _GEN_5742 : _GEN_5741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5744 = io_inputBit | _GEN_5743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5745 = i == 10'h310 ? _GEN_5744 : _GEN_5743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5746 = ~io_inputBit | _GEN_5745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5747 = i == 10'h311 ? _GEN_5746 : _GEN_5745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5748 = io_inputBit ? 1'h0 : _GEN_5747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5749 = i == 10'h311 ? _GEN_5748 : _GEN_5747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5750 = ~io_inputBit ? 1'h0 : _GEN_4753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5751 = i == 10'h1 ? _GEN_5750 : _GEN_4753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5752 = io_inputBit ? 1'h0 : _GEN_5751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5753 = i == 10'h2 ? _GEN_5752 : _GEN_5751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5754 = io_inputBit ? 1'h0 : _GEN_5753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5755 = i == 10'h5 ? _GEN_5754 : _GEN_5753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5756 = ~io_inputBit ? 1'h0 : _GEN_5755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5757 = i == 10'h9 ? _GEN_5756 : _GEN_5755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5758 = io_inputBit ? 1'h0 : _GEN_5757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5759 = i == 10'hb ? _GEN_5758 : _GEN_5757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5760 = ~io_inputBit ? 1'h0 : _GEN_5759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5761 = i == 10'h29 ? _GEN_5760 : _GEN_5759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5762 = io_inputBit ? 1'h0 : _GEN_5761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5763 = i == 10'h30 ? _GEN_5762 : _GEN_5761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5764 = ~io_inputBit ? 1'h0 : _GEN_5763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5765 = i == 10'h54 ? _GEN_5764 : _GEN_5763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5766 = io_inputBit ? 1'h0 : _GEN_5765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5767 = i == 10'h61 ? _GEN_5766 : _GEN_5765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5768 = ~io_inputBit ? 1'h0 : _GEN_5767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5769 = i == 10'haa ? _GEN_5768 : _GEN_5767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5770 = ~io_inputBit ? 1'h0 : _GEN_5769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5771 = i == 10'h156 ? _GEN_5770 : _GEN_5769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5772 = io_inputBit ? 1'h0 : _GEN_5771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5773 = i == 10'h188 ? _GEN_5772 : _GEN_5771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5774 = ~io_inputBit ? 1'h0 : _GEN_5773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5775 = i == 10'h2ae ? _GEN_5774 : _GEN_5773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5776 = io_inputBit | _GEN_5775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5777 = i == 10'h2ae ? _GEN_5776 : _GEN_5775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5778 = ~io_inputBit ? 1'h0 : _GEN_5777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5779 = i == 10'h2af ? _GEN_5778 : _GEN_5777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5780 = io_inputBit | _GEN_5779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5781 = i == 10'h2af ? _GEN_5780 : _GEN_5779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5782 = ~io_inputBit ? 1'h0 : _GEN_5781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5783 = i == 10'h2b0 ? _GEN_5782 : _GEN_5781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5784 = io_inputBit | _GEN_5783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5785 = i == 10'h2b0 ? _GEN_5784 : _GEN_5783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5786 = ~io_inputBit ? 1'h0 : _GEN_5785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5787 = i == 10'h2b1 ? _GEN_5786 : _GEN_5785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5788 = io_inputBit | _GEN_5787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5789 = i == 10'h2b1 ? _GEN_5788 : _GEN_5787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5790 = ~io_inputBit ? 1'h0 : _GEN_5789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5791 = i == 10'h2b2 ? _GEN_5790 : _GEN_5789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5792 = io_inputBit | _GEN_5791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5793 = i == 10'h2b2 ? _GEN_5792 : _GEN_5791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5794 = ~io_inputBit ? 1'h0 : _GEN_5793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5795 = i == 10'h2b3 ? _GEN_5794 : _GEN_5793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5796 = io_inputBit | _GEN_5795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5797 = i == 10'h2b3 ? _GEN_5796 : _GEN_5795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5798 = ~io_inputBit ? 1'h0 : _GEN_5797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5799 = i == 10'h2b4 ? _GEN_5798 : _GEN_5797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5800 = io_inputBit | _GEN_5799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5801 = i == 10'h2b4 ? _GEN_5800 : _GEN_5799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5802 = ~io_inputBit ? 1'h0 : _GEN_5801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5803 = i == 10'h2b5 ? _GEN_5802 : _GEN_5801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5804 = io_inputBit | _GEN_5803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5805 = i == 10'h2b5 ? _GEN_5804 : _GEN_5803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5806 = ~io_inputBit ? 1'h0 : _GEN_5805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5807 = i == 10'h2b6 ? _GEN_5806 : _GEN_5805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5808 = io_inputBit | _GEN_5807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5809 = i == 10'h2b6 ? _GEN_5808 : _GEN_5807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5810 = ~io_inputBit ? 1'h0 : _GEN_5809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5811 = i == 10'h2b7 ? _GEN_5810 : _GEN_5809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5812 = io_inputBit | _GEN_5811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5813 = i == 10'h2b7 ? _GEN_5812 : _GEN_5811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5814 = ~io_inputBit ? 1'h0 : _GEN_5813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5815 = i == 10'h2b8 ? _GEN_5814 : _GEN_5813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5816 = io_inputBit | _GEN_5815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5817 = i == 10'h2b8 ? _GEN_5816 : _GEN_5815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5818 = ~io_inputBit ? 1'h0 : _GEN_5817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5819 = i == 10'h2b9 ? _GEN_5818 : _GEN_5817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5820 = io_inputBit | _GEN_5819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5821 = i == 10'h2b9 ? _GEN_5820 : _GEN_5819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5822 = ~io_inputBit ? 1'h0 : _GEN_5821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5823 = i == 10'h2ba ? _GEN_5822 : _GEN_5821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5824 = io_inputBit | _GEN_5823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5825 = i == 10'h2ba ? _GEN_5824 : _GEN_5823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5826 = ~io_inputBit ? 1'h0 : _GEN_5825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5827 = i == 10'h2bb ? _GEN_5826 : _GEN_5825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5828 = io_inputBit | _GEN_5827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5829 = i == 10'h2bb ? _GEN_5828 : _GEN_5827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5830 = ~io_inputBit ? 1'h0 : _GEN_5829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5831 = i == 10'h2bc ? _GEN_5830 : _GEN_5829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5832 = io_inputBit | _GEN_5831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5833 = i == 10'h2bc ? _GEN_5832 : _GEN_5831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5834 = ~io_inputBit ? 1'h0 : _GEN_5833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5835 = i == 10'h2bd ? _GEN_5834 : _GEN_5833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5836 = io_inputBit | _GEN_5835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5837 = i == 10'h2bd ? _GEN_5836 : _GEN_5835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5838 = ~io_inputBit ? 1'h0 : _GEN_5837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5839 = i == 10'h2be ? _GEN_5838 : _GEN_5837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5840 = io_inputBit | _GEN_5839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5841 = i == 10'h2be ? _GEN_5840 : _GEN_5839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5842 = ~io_inputBit ? 1'h0 : _GEN_5841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5843 = i == 10'h2bf ? _GEN_5842 : _GEN_5841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5844 = io_inputBit | _GEN_5843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5845 = i == 10'h2bf ? _GEN_5844 : _GEN_5843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5846 = ~io_inputBit ? 1'h0 : _GEN_5845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5847 = i == 10'h2c0 ? _GEN_5846 : _GEN_5845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5848 = io_inputBit | _GEN_5847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5849 = i == 10'h2c0 ? _GEN_5848 : _GEN_5847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5850 = ~io_inputBit ? 1'h0 : _GEN_5849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5851 = i == 10'h2c1 ? _GEN_5850 : _GEN_5849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5852 = io_inputBit | _GEN_5851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5853 = i == 10'h2c1 ? _GEN_5852 : _GEN_5851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5854 = ~io_inputBit ? 1'h0 : _GEN_5853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5855 = i == 10'h2c2 ? _GEN_5854 : _GEN_5853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5856 = io_inputBit | _GEN_5855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5857 = i == 10'h2c2 ? _GEN_5856 : _GEN_5855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5858 = ~io_inputBit ? 1'h0 : _GEN_5857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5859 = i == 10'h2c3 ? _GEN_5858 : _GEN_5857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5860 = io_inputBit | _GEN_5859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5861 = i == 10'h2c3 ? _GEN_5860 : _GEN_5859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5862 = ~io_inputBit ? 1'h0 : _GEN_5861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5863 = i == 10'h2c4 ? _GEN_5862 : _GEN_5861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5864 = io_inputBit | _GEN_5863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5865 = i == 10'h2c4 ? _GEN_5864 : _GEN_5863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5866 = ~io_inputBit ? 1'h0 : _GEN_5865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5867 = i == 10'h2c5 ? _GEN_5866 : _GEN_5865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5868 = io_inputBit | _GEN_5867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5869 = i == 10'h2c5 ? _GEN_5868 : _GEN_5867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5870 = ~io_inputBit ? 1'h0 : _GEN_5869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5871 = i == 10'h2c6 ? _GEN_5870 : _GEN_5869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5872 = io_inputBit | _GEN_5871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5873 = i == 10'h2c6 ? _GEN_5872 : _GEN_5871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5874 = ~io_inputBit ? 1'h0 : _GEN_5873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5875 = i == 10'h2c7 ? _GEN_5874 : _GEN_5873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5876 = io_inputBit | _GEN_5875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5877 = i == 10'h2c7 ? _GEN_5876 : _GEN_5875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5878 = ~io_inputBit ? 1'h0 : _GEN_5877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5879 = i == 10'h2c8 ? _GEN_5878 : _GEN_5877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5880 = io_inputBit | _GEN_5879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5881 = i == 10'h2c8 ? _GEN_5880 : _GEN_5879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5882 = ~io_inputBit ? 1'h0 : _GEN_5881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5883 = i == 10'h2c9 ? _GEN_5882 : _GEN_5881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5884 = io_inputBit | _GEN_5883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5885 = i == 10'h2c9 ? _GEN_5884 : _GEN_5883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5886 = ~io_inputBit ? 1'h0 : _GEN_5885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5887 = i == 10'h2ca ? _GEN_5886 : _GEN_5885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5888 = io_inputBit | _GEN_5887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5889 = i == 10'h2ca ? _GEN_5888 : _GEN_5887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5890 = ~io_inputBit ? 1'h0 : _GEN_5889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5891 = i == 10'h2cb ? _GEN_5890 : _GEN_5889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5892 = io_inputBit | _GEN_5891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5893 = i == 10'h2cb ? _GEN_5892 : _GEN_5891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5894 = ~io_inputBit ? 1'h0 : _GEN_5893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5895 = i == 10'h2cc ? _GEN_5894 : _GEN_5893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5896 = io_inputBit | _GEN_5895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5897 = i == 10'h2cc ? _GEN_5896 : _GEN_5895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5898 = ~io_inputBit ? 1'h0 : _GEN_5897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5899 = i == 10'h2cd ? _GEN_5898 : _GEN_5897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5900 = io_inputBit | _GEN_5899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5901 = i == 10'h2cd ? _GEN_5900 : _GEN_5899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5902 = ~io_inputBit ? 1'h0 : _GEN_5901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5903 = i == 10'h2ce ? _GEN_5902 : _GEN_5901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5904 = io_inputBit | _GEN_5903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5905 = i == 10'h2ce ? _GEN_5904 : _GEN_5903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5906 = ~io_inputBit ? 1'h0 : _GEN_5905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5907 = i == 10'h2cf ? _GEN_5906 : _GEN_5905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5908 = io_inputBit | _GEN_5907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5909 = i == 10'h2cf ? _GEN_5908 : _GEN_5907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5910 = ~io_inputBit ? 1'h0 : _GEN_5909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5911 = i == 10'h2d0 ? _GEN_5910 : _GEN_5909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5912 = io_inputBit | _GEN_5911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5913 = i == 10'h2d0 ? _GEN_5912 : _GEN_5911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5914 = ~io_inputBit ? 1'h0 : _GEN_5913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5915 = i == 10'h2d1 ? _GEN_5914 : _GEN_5913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5916 = io_inputBit | _GEN_5915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5917 = i == 10'h2d1 ? _GEN_5916 : _GEN_5915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5918 = ~io_inputBit ? 1'h0 : _GEN_5917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5919 = i == 10'h2d2 ? _GEN_5918 : _GEN_5917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5920 = io_inputBit | _GEN_5919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5921 = i == 10'h2d2 ? _GEN_5920 : _GEN_5919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5922 = ~io_inputBit ? 1'h0 : _GEN_5921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5923 = i == 10'h2d3 ? _GEN_5922 : _GEN_5921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5924 = io_inputBit | _GEN_5923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5925 = i == 10'h2d3 ? _GEN_5924 : _GEN_5923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5926 = ~io_inputBit ? 1'h0 : _GEN_5925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5927 = i == 10'h2d4 ? _GEN_5926 : _GEN_5925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5928 = io_inputBit | _GEN_5927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5929 = i == 10'h2d4 ? _GEN_5928 : _GEN_5927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5930 = ~io_inputBit ? 1'h0 : _GEN_5929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5931 = i == 10'h2d5 ? _GEN_5930 : _GEN_5929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5932 = io_inputBit | _GEN_5931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5933 = i == 10'h2d5 ? _GEN_5932 : _GEN_5931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5934 = ~io_inputBit ? 1'h0 : _GEN_5933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5935 = i == 10'h2d6 ? _GEN_5934 : _GEN_5933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5936 = io_inputBit | _GEN_5935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5937 = i == 10'h2d6 ? _GEN_5936 : _GEN_5935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5938 = ~io_inputBit ? 1'h0 : _GEN_5937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5939 = i == 10'h2d7 ? _GEN_5938 : _GEN_5937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5940 = io_inputBit | _GEN_5939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5941 = i == 10'h2d7 ? _GEN_5940 : _GEN_5939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5942 = ~io_inputBit ? 1'h0 : _GEN_5941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5943 = i == 10'h2d8 ? _GEN_5942 : _GEN_5941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5944 = io_inputBit | _GEN_5943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5945 = i == 10'h2d8 ? _GEN_5944 : _GEN_5943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5946 = ~io_inputBit ? 1'h0 : _GEN_5945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5947 = i == 10'h2d9 ? _GEN_5946 : _GEN_5945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5948 = io_inputBit | _GEN_5947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5949 = i == 10'h2d9 ? _GEN_5948 : _GEN_5947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5950 = ~io_inputBit ? 1'h0 : _GEN_5949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5951 = i == 10'h2da ? _GEN_5950 : _GEN_5949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5952 = io_inputBit | _GEN_5951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5953 = i == 10'h2da ? _GEN_5952 : _GEN_5951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5954 = ~io_inputBit ? 1'h0 : _GEN_5953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5955 = i == 10'h2db ? _GEN_5954 : _GEN_5953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5956 = io_inputBit | _GEN_5955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5957 = i == 10'h2db ? _GEN_5956 : _GEN_5955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5958 = ~io_inputBit ? 1'h0 : _GEN_5957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5959 = i == 10'h2dc ? _GEN_5958 : _GEN_5957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5960 = io_inputBit | _GEN_5959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5961 = i == 10'h2dc ? _GEN_5960 : _GEN_5959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5962 = ~io_inputBit ? 1'h0 : _GEN_5961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5963 = i == 10'h2dd ? _GEN_5962 : _GEN_5961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5964 = io_inputBit | _GEN_5963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5965 = i == 10'h2dd ? _GEN_5964 : _GEN_5963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5966 = ~io_inputBit ? 1'h0 : _GEN_5965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5967 = i == 10'h2de ? _GEN_5966 : _GEN_5965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5968 = io_inputBit | _GEN_5967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5969 = i == 10'h2de ? _GEN_5968 : _GEN_5967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5970 = ~io_inputBit ? 1'h0 : _GEN_5969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5971 = i == 10'h2df ? _GEN_5970 : _GEN_5969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5972 = io_inputBit | _GEN_5971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5973 = i == 10'h2df ? _GEN_5972 : _GEN_5971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5974 = ~io_inputBit ? 1'h0 : _GEN_5973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5975 = i == 10'h2e0 ? _GEN_5974 : _GEN_5973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5976 = io_inputBit | _GEN_5975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5977 = i == 10'h2e0 ? _GEN_5976 : _GEN_5975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5978 = ~io_inputBit ? 1'h0 : _GEN_5977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5979 = i == 10'h2e1 ? _GEN_5978 : _GEN_5977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5980 = io_inputBit | _GEN_5979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5981 = i == 10'h2e1 ? _GEN_5980 : _GEN_5979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5982 = ~io_inputBit ? 1'h0 : _GEN_5981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5983 = i == 10'h2e2 ? _GEN_5982 : _GEN_5981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5984 = io_inputBit | _GEN_5983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5985 = i == 10'h2e2 ? _GEN_5984 : _GEN_5983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5986 = ~io_inputBit ? 1'h0 : _GEN_5985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5987 = i == 10'h2e3 ? _GEN_5986 : _GEN_5985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5988 = io_inputBit | _GEN_5987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5989 = i == 10'h2e3 ? _GEN_5988 : _GEN_5987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5990 = ~io_inputBit ? 1'h0 : _GEN_5989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5991 = i == 10'h2e4 ? _GEN_5990 : _GEN_5989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5992 = io_inputBit | _GEN_5991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5993 = i == 10'h2e4 ? _GEN_5992 : _GEN_5991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5994 = ~io_inputBit ? 1'h0 : _GEN_5993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5995 = i == 10'h2e5 ? _GEN_5994 : _GEN_5993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5996 = io_inputBit | _GEN_5995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5997 = i == 10'h2e5 ? _GEN_5996 : _GEN_5995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_5998 = ~io_inputBit ? 1'h0 : _GEN_5997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5999 = i == 10'h2e6 ? _GEN_5998 : _GEN_5997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6000 = io_inputBit | _GEN_5999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6001 = i == 10'h2e6 ? _GEN_6000 : _GEN_5999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6002 = ~io_inputBit ? 1'h0 : _GEN_6001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6003 = i == 10'h2e7 ? _GEN_6002 : _GEN_6001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6004 = io_inputBit | _GEN_6003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6005 = i == 10'h2e7 ? _GEN_6004 : _GEN_6003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6006 = ~io_inputBit ? 1'h0 : _GEN_6005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6007 = i == 10'h2e8 ? _GEN_6006 : _GEN_6005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6008 = io_inputBit | _GEN_6007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6009 = i == 10'h2e8 ? _GEN_6008 : _GEN_6007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6010 = ~io_inputBit ? 1'h0 : _GEN_6009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6011 = i == 10'h2e9 ? _GEN_6010 : _GEN_6009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6012 = io_inputBit | _GEN_6011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6013 = i == 10'h2e9 ? _GEN_6012 : _GEN_6011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6014 = ~io_inputBit ? 1'h0 : _GEN_6013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6015 = i == 10'h2ea ? _GEN_6014 : _GEN_6013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6016 = io_inputBit | _GEN_6015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6017 = i == 10'h2ea ? _GEN_6016 : _GEN_6015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6018 = ~io_inputBit ? 1'h0 : _GEN_6017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6019 = i == 10'h2eb ? _GEN_6018 : _GEN_6017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6020 = io_inputBit | _GEN_6019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6021 = i == 10'h2eb ? _GEN_6020 : _GEN_6019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6022 = ~io_inputBit ? 1'h0 : _GEN_6021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6023 = i == 10'h2ec ? _GEN_6022 : _GEN_6021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6024 = io_inputBit | _GEN_6023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6025 = i == 10'h2ec ? _GEN_6024 : _GEN_6023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6026 = ~io_inputBit ? 1'h0 : _GEN_6025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6027 = i == 10'h2ed ? _GEN_6026 : _GEN_6025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6028 = io_inputBit | _GEN_6027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6029 = i == 10'h2ed ? _GEN_6028 : _GEN_6027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6030 = ~io_inputBit ? 1'h0 : _GEN_6029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6031 = i == 10'h2ee ? _GEN_6030 : _GEN_6029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6032 = io_inputBit | _GEN_6031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6033 = i == 10'h2ee ? _GEN_6032 : _GEN_6031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6034 = ~io_inputBit ? 1'h0 : _GEN_6033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6035 = i == 10'h2ef ? _GEN_6034 : _GEN_6033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6036 = io_inputBit | _GEN_6035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6037 = i == 10'h2ef ? _GEN_6036 : _GEN_6035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6038 = ~io_inputBit ? 1'h0 : _GEN_6037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6039 = i == 10'h2f0 ? _GEN_6038 : _GEN_6037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6040 = io_inputBit | _GEN_6039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6041 = i == 10'h2f0 ? _GEN_6040 : _GEN_6039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6042 = ~io_inputBit ? 1'h0 : _GEN_6041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6043 = i == 10'h2f1 ? _GEN_6042 : _GEN_6041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6044 = io_inputBit | _GEN_6043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6045 = i == 10'h2f1 ? _GEN_6044 : _GEN_6043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6046 = ~io_inputBit ? 1'h0 : _GEN_6045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6047 = i == 10'h2f2 ? _GEN_6046 : _GEN_6045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6048 = io_inputBit | _GEN_6047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6049 = i == 10'h2f2 ? _GEN_6048 : _GEN_6047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6050 = ~io_inputBit ? 1'h0 : _GEN_6049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6051 = i == 10'h2f3 ? _GEN_6050 : _GEN_6049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6052 = io_inputBit | _GEN_6051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6053 = i == 10'h2f3 ? _GEN_6052 : _GEN_6051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6054 = ~io_inputBit ? 1'h0 : _GEN_6053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6055 = i == 10'h2f4 ? _GEN_6054 : _GEN_6053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6056 = io_inputBit | _GEN_6055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6057 = i == 10'h2f4 ? _GEN_6056 : _GEN_6055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6058 = ~io_inputBit ? 1'h0 : _GEN_6057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6059 = i == 10'h2f5 ? _GEN_6058 : _GEN_6057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6060 = io_inputBit | _GEN_6059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6061 = i == 10'h2f5 ? _GEN_6060 : _GEN_6059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6062 = ~io_inputBit ? 1'h0 : _GEN_6061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6063 = i == 10'h2f6 ? _GEN_6062 : _GEN_6061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6064 = io_inputBit | _GEN_6063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6065 = i == 10'h2f6 ? _GEN_6064 : _GEN_6063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6066 = ~io_inputBit ? 1'h0 : _GEN_6065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6067 = i == 10'h2f7 ? _GEN_6066 : _GEN_6065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6068 = io_inputBit | _GEN_6067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6069 = i == 10'h2f7 ? _GEN_6068 : _GEN_6067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6070 = ~io_inputBit ? 1'h0 : _GEN_6069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6071 = i == 10'h2f8 ? _GEN_6070 : _GEN_6069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6072 = io_inputBit | _GEN_6071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6073 = i == 10'h2f8 ? _GEN_6072 : _GEN_6071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6074 = ~io_inputBit ? 1'h0 : _GEN_6073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6075 = i == 10'h2f9 ? _GEN_6074 : _GEN_6073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6076 = io_inputBit | _GEN_6075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6077 = i == 10'h2f9 ? _GEN_6076 : _GEN_6075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6078 = ~io_inputBit ? 1'h0 : _GEN_6077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6079 = i == 10'h2fa ? _GEN_6078 : _GEN_6077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6080 = io_inputBit | _GEN_6079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6081 = i == 10'h2fa ? _GEN_6080 : _GEN_6079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6082 = ~io_inputBit ? 1'h0 : _GEN_6081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6083 = i == 10'h2fb ? _GEN_6082 : _GEN_6081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6084 = io_inputBit | _GEN_6083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6085 = i == 10'h2fb ? _GEN_6084 : _GEN_6083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6086 = ~io_inputBit ? 1'h0 : _GEN_6085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6087 = i == 10'h2fc ? _GEN_6086 : _GEN_6085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6088 = io_inputBit | _GEN_6087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6089 = i == 10'h2fc ? _GEN_6088 : _GEN_6087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6090 = ~io_inputBit ? 1'h0 : _GEN_6089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6091 = i == 10'h2fd ? _GEN_6090 : _GEN_6089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6092 = io_inputBit | _GEN_6091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6093 = i == 10'h2fd ? _GEN_6092 : _GEN_6091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6094 = ~io_inputBit ? 1'h0 : _GEN_6093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6095 = i == 10'h2fe ? _GEN_6094 : _GEN_6093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6096 = io_inputBit | _GEN_6095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6097 = i == 10'h2fe ? _GEN_6096 : _GEN_6095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6098 = ~io_inputBit ? 1'h0 : _GEN_6097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6099 = i == 10'h2ff ? _GEN_6098 : _GEN_6097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6100 = io_inputBit | _GEN_6099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6101 = i == 10'h2ff ? _GEN_6100 : _GEN_6099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6102 = ~io_inputBit ? 1'h0 : _GEN_6101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6103 = i == 10'h300 ? _GEN_6102 : _GEN_6101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6104 = io_inputBit | _GEN_6103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6105 = i == 10'h300 ? _GEN_6104 : _GEN_6103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6106 = ~io_inputBit ? 1'h0 : _GEN_6105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6107 = i == 10'h301 ? _GEN_6106 : _GEN_6105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6108 = io_inputBit | _GEN_6107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6109 = i == 10'h301 ? _GEN_6108 : _GEN_6107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6110 = ~io_inputBit ? 1'h0 : _GEN_6109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6111 = i == 10'h302 ? _GEN_6110 : _GEN_6109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6112 = io_inputBit | _GEN_6111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6113 = i == 10'h302 ? _GEN_6112 : _GEN_6111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6114 = ~io_inputBit ? 1'h0 : _GEN_6113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6115 = i == 10'h303 ? _GEN_6114 : _GEN_6113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6116 = io_inputBit | _GEN_6115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6117 = i == 10'h303 ? _GEN_6116 : _GEN_6115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6118 = ~io_inputBit ? 1'h0 : _GEN_6117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6119 = i == 10'h304 ? _GEN_6118 : _GEN_6117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6120 = io_inputBit | _GEN_6119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6121 = i == 10'h304 ? _GEN_6120 : _GEN_6119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6122 = ~io_inputBit ? 1'h0 : _GEN_6121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6123 = i == 10'h305 ? _GEN_6122 : _GEN_6121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6124 = io_inputBit | _GEN_6123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6125 = i == 10'h305 ? _GEN_6124 : _GEN_6123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6126 = ~io_inputBit ? 1'h0 : _GEN_6125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6127 = i == 10'h306 ? _GEN_6126 : _GEN_6125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6128 = io_inputBit | _GEN_6127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6129 = i == 10'h306 ? _GEN_6128 : _GEN_6127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6130 = ~io_inputBit ? 1'h0 : _GEN_6129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6131 = i == 10'h307 ? _GEN_6130 : _GEN_6129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6132 = io_inputBit | _GEN_6131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6133 = i == 10'h307 ? _GEN_6132 : _GEN_6131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6134 = ~io_inputBit ? 1'h0 : _GEN_6133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6135 = i == 10'h308 ? _GEN_6134 : _GEN_6133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6136 = io_inputBit | _GEN_6135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6137 = i == 10'h308 ? _GEN_6136 : _GEN_6135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6138 = ~io_inputBit ? 1'h0 : _GEN_6137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6139 = i == 10'h309 ? _GEN_6138 : _GEN_6137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6140 = io_inputBit | _GEN_6139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6141 = i == 10'h309 ? _GEN_6140 : _GEN_6139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6142 = ~io_inputBit ? 1'h0 : _GEN_6141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6143 = i == 10'h30a ? _GEN_6142 : _GEN_6141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6144 = io_inputBit | _GEN_6143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6145 = i == 10'h30a ? _GEN_6144 : _GEN_6143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6146 = ~io_inputBit ? 1'h0 : _GEN_6145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6147 = i == 10'h30b ? _GEN_6146 : _GEN_6145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6148 = io_inputBit | _GEN_6147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6149 = i == 10'h30b ? _GEN_6148 : _GEN_6147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6150 = ~io_inputBit ? 1'h0 : _GEN_6149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6151 = i == 10'h30c ? _GEN_6150 : _GEN_6149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6152 = io_inputBit | _GEN_6151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6153 = i == 10'h30c ? _GEN_6152 : _GEN_6151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6154 = ~io_inputBit ? 1'h0 : _GEN_6153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6155 = i == 10'h30d ? _GEN_6154 : _GEN_6153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6156 = io_inputBit | _GEN_6155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6157 = i == 10'h30d ? _GEN_6156 : _GEN_6155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6158 = ~io_inputBit ? 1'h0 : _GEN_6157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6159 = i == 10'h30e ? _GEN_6158 : _GEN_6157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6160 = io_inputBit | _GEN_6159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6161 = i == 10'h30e ? _GEN_6160 : _GEN_6159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6162 = ~io_inputBit ? 1'h0 : _GEN_6161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6163 = i == 10'h30f ? _GEN_6162 : _GEN_6161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6164 = io_inputBit | _GEN_6163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6165 = i == 10'h30f ? _GEN_6164 : _GEN_6163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6166 = ~io_inputBit ? 1'h0 : _GEN_6165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6167 = i == 10'h310 ? _GEN_6166 : _GEN_6165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6168 = io_inputBit | _GEN_6167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6169 = i == 10'h310 ? _GEN_6168 : _GEN_6167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6170 = ~io_inputBit ? 1'h0 : _GEN_6169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6171 = i == 10'h311 ? _GEN_6170 : _GEN_6169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6172 = io_inputBit | _GEN_6171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6173 = i == 10'h311 ? _GEN_6172 : _GEN_6171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6174 = ~io_inputBit ? 1'h0 : _GEN_4785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6175 = i == 10'h0 ? _GEN_6174 : _GEN_4785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6176 = io_inputBit | _GEN_6175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6177 = i == 10'h2 ? _GEN_6176 : _GEN_6175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6178 = io_inputBit | _GEN_6177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6179 = i == 10'h5 ? _GEN_6178 : _GEN_6177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6180 = io_inputBit | _GEN_6179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6181 = i == 10'hb ? _GEN_6180 : _GEN_6179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6182 = ~io_inputBit ? 1'h0 : _GEN_6181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6183 = i == 10'h17 ? _GEN_6182 : _GEN_6181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6184 = ~io_inputBit ? 1'h0 : _GEN_6183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6185 = i == 10'h30 ? _GEN_6184 : _GEN_6183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6186 = io_inputBit | _GEN_6185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6187 = i == 10'h62 ? _GEN_6186 : _GEN_6185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6188 = ~io_inputBit ? 1'h0 : _GEN_6187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6189 = i == 10'hc5 ? _GEN_6188 : _GEN_6187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6190 = io_inputBit | _GEN_6189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6192 = ~io_inputBit ? 1'h0 : _GEN_4865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6193 = i == 10'h0 ? _GEN_6192 : _GEN_4865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6194 = io_inputBit | _GEN_6193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6195 = i == 10'h2 ? _GEN_6194 : _GEN_6193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6196 = io_inputBit | _GEN_6195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6197 = i == 10'h5 ? _GEN_6196 : _GEN_6195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6198 = io_inputBit | _GEN_6197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6199 = i == 10'h18 ? _GEN_6198 : _GEN_6197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6200 = ~io_inputBit ? 1'h0 : _GEN_6199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6201 = i == 10'h2f ? _GEN_6200 : _GEN_6199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6202 = ~io_inputBit | _GEN_6201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6203 = i == 10'h30 ? _GEN_6202 : _GEN_6201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6204 = ~io_inputBit ? 1'h0 : _GEN_6203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6205 = i == 10'h31 ? _GEN_6204 : _GEN_6203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6206 = io_inputBit | _GEN_6205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6207 = i == 10'h60 ? _GEN_6206 : _GEN_6205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6208 = io_inputBit ? 1'h0 : _GEN_6207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6209 = i == 10'h62 ? _GEN_6208 : _GEN_6207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6210 = io_inputBit | _GEN_6209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6211 = i == 10'h64 ? _GEN_6210 : _GEN_6209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6212 = ~io_inputBit ? 1'h0 : _GEN_6211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6213 = i == 10'hc1 ? _GEN_6212 : _GEN_6211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6214 = io_inputBit | _GEN_6213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6215 = i == 10'hc1 ? _GEN_6214 : _GEN_6213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6216 = ~io_inputBit | _GEN_6215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6217 = i == 10'hc5 ? _GEN_6216 : _GEN_6215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6218 = io_inputBit ? 1'h0 : _GEN_6217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6219 = i == 10'hc5 ? _GEN_6218 : _GEN_6217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6220 = ~io_inputBit ? 1'h0 : _GEN_6219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6221 = i == 10'hc9 ? _GEN_6220 : _GEN_6219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6222 = io_inputBit | _GEN_6221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6224 = ~io_inputBit ? 1'h0 : _GEN_4987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6225 = i == 10'h0 ? _GEN_6224 : _GEN_4987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6226 = io_inputBit ? 1'h0 : _GEN_6225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6227 = i == 10'h2 ? _GEN_6226 : _GEN_6225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6228 = io_inputBit ? 1'h0 : _GEN_6227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6229 = i == 10'h5 ? _GEN_6228 : _GEN_6227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6230 = io_inputBit ? 1'h0 : _GEN_6229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6231 = i == 10'h18 ? _GEN_6230 : _GEN_6229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6232 = io_inputBit | _GEN_6231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6233 = i == 10'h5f ? _GEN_6232 : _GEN_6231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6234 = io_inputBit ? 1'h0 : _GEN_6233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6235 = i == 10'h60 ? _GEN_6234 : _GEN_6233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6236 = io_inputBit | _GEN_6235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6237 = i == 10'h61 ? _GEN_6236 : _GEN_6235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6238 = io_inputBit ? 1'h0 : _GEN_6237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6239 = i == 10'h62 ? _GEN_6238 : _GEN_6237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6240 = io_inputBit | _GEN_6239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6241 = i == 10'h63 ? _GEN_6240 : _GEN_6239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6242 = io_inputBit ? 1'h0 : _GEN_6241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6243 = i == 10'h64 ? _GEN_6242 : _GEN_6241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6244 = ~io_inputBit ? 1'h0 : _GEN_6243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6245 = i == 10'hbf ? _GEN_6244 : _GEN_6243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6246 = io_inputBit | _GEN_6245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6247 = i == 10'hbf ? _GEN_6246 : _GEN_6245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6248 = ~io_inputBit | _GEN_6247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6249 = i == 10'hc1 ? _GEN_6248 : _GEN_6247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6250 = io_inputBit ? 1'h0 : _GEN_6249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6251 = i == 10'hc1 ? _GEN_6250 : _GEN_6249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6252 = ~io_inputBit ? 1'h0 : _GEN_6251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6253 = i == 10'hc3 ? _GEN_6252 : _GEN_6251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6254 = io_inputBit | _GEN_6253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6255 = i == 10'hc3 ? _GEN_6254 : _GEN_6253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6256 = ~io_inputBit | _GEN_6255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6257 = i == 10'hc5 ? _GEN_6256 : _GEN_6255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6258 = io_inputBit ? 1'h0 : _GEN_6257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6259 = i == 10'hc5 ? _GEN_6258 : _GEN_6257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6260 = ~io_inputBit ? 1'h0 : _GEN_6259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6261 = i == 10'hc7 ? _GEN_6260 : _GEN_6259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6262 = io_inputBit | _GEN_6261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6263 = i == 10'hc7 ? _GEN_6262 : _GEN_6261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6264 = ~io_inputBit | _GEN_6263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6265 = i == 10'hc9 ? _GEN_6264 : _GEN_6263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6268 = ~io_inputBit ? 1'h0 : _GEN_5169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6269 = i == 10'h1 ? _GEN_6268 : _GEN_5169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6270 = io_inputBit ? 1'h0 : _GEN_6269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6271 = i == 10'h2 ? _GEN_6270 : _GEN_6269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6272 = ~io_inputBit ? 1'h0 : _GEN_6271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6273 = i == 10'h4 ? _GEN_6272 : _GEN_6271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6274 = io_inputBit ? 1'h0 : _GEN_6273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6275 = i == 10'h5 ? _GEN_6274 : _GEN_6273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6276 = ~io_inputBit ? 1'h0 : _GEN_6275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6277 = i == 10'ha ? _GEN_6276 : _GEN_6275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6278 = ~io_inputBit ? 1'h0 : _GEN_6277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6279 = i == 10'h16 ? _GEN_6278 : _GEN_6277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6280 = io_inputBit ? 1'h0 : _GEN_6279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6281 = i == 10'h18 ? _GEN_6280 : _GEN_6279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6282 = ~io_inputBit ? 1'h0 : _GEN_6281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6283 = i == 10'h2e ? _GEN_6282 : _GEN_6281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6284 = ~io_inputBit ? 1'h0 : _GEN_6283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6285 = i == 10'h5e ? _GEN_6284 : _GEN_6283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6286 = io_inputBit ? 1'h0 : _GEN_6285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6287 = i == 10'h64 ? _GEN_6286 : _GEN_6285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6288 = ~io_inputBit ? 1'h0 : _GEN_6287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6289 = i == 10'hbe ? _GEN_6288 : _GEN_6287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6290 = io_inputBit | _GEN_6289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6291 = i == 10'hbe ? _GEN_6290 : _GEN_6289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6292 = ~io_inputBit | _GEN_6291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6293 = i == 10'hbf ? _GEN_6292 : _GEN_6291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6294 = io_inputBit ? 1'h0 : _GEN_6293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6295 = i == 10'hbf ? _GEN_6294 : _GEN_6293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6296 = ~io_inputBit ? 1'h0 : _GEN_6295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6297 = i == 10'hc0 ? _GEN_6296 : _GEN_6295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6298 = io_inputBit | _GEN_6297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6299 = i == 10'hc0 ? _GEN_6298 : _GEN_6297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6300 = ~io_inputBit | _GEN_6299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6301 = i == 10'hc1 ? _GEN_6300 : _GEN_6299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6302 = io_inputBit ? 1'h0 : _GEN_6301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6303 = i == 10'hc1 ? _GEN_6302 : _GEN_6301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6304 = ~io_inputBit ? 1'h0 : _GEN_6303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6305 = i == 10'hc2 ? _GEN_6304 : _GEN_6303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6306 = io_inputBit | _GEN_6305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6307 = i == 10'hc2 ? _GEN_6306 : _GEN_6305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6308 = ~io_inputBit | _GEN_6307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6309 = i == 10'hc3 ? _GEN_6308 : _GEN_6307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6310 = io_inputBit ? 1'h0 : _GEN_6309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6311 = i == 10'hc3 ? _GEN_6310 : _GEN_6309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6312 = ~io_inputBit ? 1'h0 : _GEN_6311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6313 = i == 10'hc4 ? _GEN_6312 : _GEN_6311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6314 = io_inputBit | _GEN_6313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6315 = i == 10'hc4 ? _GEN_6314 : _GEN_6313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6316 = ~io_inputBit | _GEN_6315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6317 = i == 10'hc5 ? _GEN_6316 : _GEN_6315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6318 = io_inputBit ? 1'h0 : _GEN_6317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6319 = i == 10'hc5 ? _GEN_6318 : _GEN_6317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6320 = ~io_inputBit ? 1'h0 : _GEN_6319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6321 = i == 10'hc6 ? _GEN_6320 : _GEN_6319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6322 = io_inputBit | _GEN_6321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6323 = i == 10'hc6 ? _GEN_6322 : _GEN_6321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6324 = ~io_inputBit | _GEN_6323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6325 = i == 10'hc7 ? _GEN_6324 : _GEN_6323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6326 = io_inputBit ? 1'h0 : _GEN_6325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6327 = i == 10'hc7 ? _GEN_6326 : _GEN_6325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6328 = ~io_inputBit ? 1'h0 : _GEN_6327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6329 = i == 10'hc8 ? _GEN_6328 : _GEN_6327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6330 = io_inputBit | _GEN_6329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6331 = i == 10'hc8 ? _GEN_6330 : _GEN_6329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6332 = ~io_inputBit | _GEN_6331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6333 = i == 10'hc9 ? _GEN_6332 : _GEN_6331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6336 = ~io_inputBit ? 1'h0 : _GEN_5433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6337 = i == 10'h1 ? _GEN_6336 : _GEN_5433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6338 = io_inputBit | _GEN_6337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6339 = i == 10'h2 ? _GEN_6338 : _GEN_6337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6340 = ~io_inputBit ? 1'h0 : _GEN_6339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6341 = i == 10'h4 ? _GEN_6340 : _GEN_6339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6342 = io_inputBit | _GEN_6341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6343 = i == 10'h5 ? _GEN_6342 : _GEN_6341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6344 = ~io_inputBit ? 1'h0 : _GEN_6343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6345 = i == 10'ha ? _GEN_6344 : _GEN_6343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6346 = ~io_inputBit ? 1'h0 : _GEN_6345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6347 = i == 10'h16 ? _GEN_6346 : _GEN_6345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6348 = io_inputBit | _GEN_6347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6349 = i == 10'h18 ? _GEN_6348 : _GEN_6347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6350 = ~io_inputBit ? 1'h0 : _GEN_6349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6351 = i == 10'h2e ? _GEN_6350 : _GEN_6349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6352 = ~io_inputBit ? 1'h0 : _GEN_6351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6353 = i == 10'h5e ? _GEN_6352 : _GEN_6351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6354 = io_inputBit | _GEN_6353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6355 = i == 10'h64 ? _GEN_6354 : _GEN_6353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6356 = ~io_inputBit | _GEN_6355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6357 = i == 10'hbe ? _GEN_6356 : _GEN_6355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6358 = io_inputBit ? 1'h0 : _GEN_6357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6359 = i == 10'hbe ? _GEN_6358 : _GEN_6357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6360 = ~io_inputBit | _GEN_6359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6361 = i == 10'hbf ? _GEN_6360 : _GEN_6359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6362 = io_inputBit ? 1'h0 : _GEN_6361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6363 = i == 10'hbf ? _GEN_6362 : _GEN_6361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6364 = ~io_inputBit | _GEN_6363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6365 = i == 10'hc0 ? _GEN_6364 : _GEN_6363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6366 = io_inputBit ? 1'h0 : _GEN_6365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6367 = i == 10'hc0 ? _GEN_6366 : _GEN_6365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6368 = ~io_inputBit | _GEN_6367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6369 = i == 10'hc1 ? _GEN_6368 : _GEN_6367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6370 = io_inputBit ? 1'h0 : _GEN_6369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6371 = i == 10'hc1 ? _GEN_6370 : _GEN_6369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6372 = ~io_inputBit | _GEN_6371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6373 = i == 10'hc2 ? _GEN_6372 : _GEN_6371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6374 = io_inputBit ? 1'h0 : _GEN_6373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6375 = i == 10'hc2 ? _GEN_6374 : _GEN_6373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6376 = ~io_inputBit | _GEN_6375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6377 = i == 10'hc3 ? _GEN_6376 : _GEN_6375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6378 = io_inputBit ? 1'h0 : _GEN_6377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6379 = i == 10'hc3 ? _GEN_6378 : _GEN_6377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6380 = ~io_inputBit | _GEN_6379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6381 = i == 10'hc4 ? _GEN_6380 : _GEN_6379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6382 = io_inputBit ? 1'h0 : _GEN_6381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6383 = i == 10'hc4 ? _GEN_6382 : _GEN_6381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6384 = ~io_inputBit | _GEN_6383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6385 = i == 10'hc5 ? _GEN_6384 : _GEN_6383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6386 = io_inputBit ? 1'h0 : _GEN_6385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6387 = i == 10'hc5 ? _GEN_6386 : _GEN_6385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6388 = ~io_inputBit | _GEN_6387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6389 = i == 10'hc6 ? _GEN_6388 : _GEN_6387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6390 = io_inputBit ? 1'h0 : _GEN_6389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6391 = i == 10'hc6 ? _GEN_6390 : _GEN_6389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6392 = ~io_inputBit | _GEN_6391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6393 = i == 10'hc7 ? _GEN_6392 : _GEN_6391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6394 = io_inputBit ? 1'h0 : _GEN_6393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6395 = i == 10'hc7 ? _GEN_6394 : _GEN_6393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6396 = ~io_inputBit | _GEN_6395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6397 = i == 10'hc8 ? _GEN_6396 : _GEN_6395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6398 = io_inputBit ? 1'h0 : _GEN_6397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6399 = i == 10'hc8 ? _GEN_6398 : _GEN_6397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6400 = ~io_inputBit | _GEN_6399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6401 = i == 10'hc9 ? _GEN_6400 : _GEN_6399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6404 = ~io_inputBit ? 1'h0 : _GEN_5749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6405 = i == 10'h1 ? _GEN_6404 : _GEN_5749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6406 = io_inputBit ? 1'h0 : _GEN_6405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6407 = i == 10'h2 ? _GEN_6406 : _GEN_6405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6408 = ~io_inputBit ? 1'h0 : _GEN_6407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6409 = i == 10'h4 ? _GEN_6408 : _GEN_6407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6410 = io_inputBit ? 1'h0 : _GEN_6409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6411 = i == 10'h5 ? _GEN_6410 : _GEN_6409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6412 = ~io_inputBit ? 1'h0 : _GEN_6411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6413 = i == 10'ha ? _GEN_6412 : _GEN_6411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6414 = ~io_inputBit ? 1'h0 : _GEN_6413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6415 = i == 10'h16 ? _GEN_6414 : _GEN_6413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6416 = io_inputBit ? 1'h0 : _GEN_6415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6417 = i == 10'h18 ? _GEN_6416 : _GEN_6415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6418 = ~io_inputBit ? 1'h0 : _GEN_6417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6419 = i == 10'h2e ? _GEN_6418 : _GEN_6417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6420 = io_inputBit ? 1'h0 : _GEN_6419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6421 = i == 10'h64 ? _GEN_6420 : _GEN_6419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6422 = ~io_inputBit ? 1'h0 : _GEN_6421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6423 = i == 10'hbd ? _GEN_6422 : _GEN_6421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6424 = ~io_inputBit ? 1'h0 : _GEN_6423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6425 = i == 10'h17c ? _GEN_6424 : _GEN_6423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6426 = io_inputBit | _GEN_6425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6427 = i == 10'h17c ? _GEN_6426 : _GEN_6425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6428 = ~io_inputBit ? 1'h0 : _GEN_6427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6429 = i == 10'h17d ? _GEN_6428 : _GEN_6427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6430 = io_inputBit | _GEN_6429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6431 = i == 10'h17d ? _GEN_6430 : _GEN_6429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6432 = ~io_inputBit ? 1'h0 : _GEN_6431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6433 = i == 10'h17e ? _GEN_6432 : _GEN_6431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6434 = io_inputBit | _GEN_6433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6435 = i == 10'h17e ? _GEN_6434 : _GEN_6433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6436 = ~io_inputBit ? 1'h0 : _GEN_6435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6437 = i == 10'h17f ? _GEN_6436 : _GEN_6435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6438 = io_inputBit | _GEN_6437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6439 = i == 10'h17f ? _GEN_6438 : _GEN_6437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6440 = ~io_inputBit ? 1'h0 : _GEN_6439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6441 = i == 10'h180 ? _GEN_6440 : _GEN_6439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6442 = io_inputBit | _GEN_6441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6443 = i == 10'h180 ? _GEN_6442 : _GEN_6441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6444 = ~io_inputBit ? 1'h0 : _GEN_6443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6445 = i == 10'h181 ? _GEN_6444 : _GEN_6443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6446 = io_inputBit | _GEN_6445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6447 = i == 10'h181 ? _GEN_6446 : _GEN_6445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6448 = ~io_inputBit ? 1'h0 : _GEN_6447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6449 = i == 10'h182 ? _GEN_6448 : _GEN_6447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6450 = io_inputBit | _GEN_6449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6451 = i == 10'h182 ? _GEN_6450 : _GEN_6449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6452 = ~io_inputBit ? 1'h0 : _GEN_6451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6453 = i == 10'h183 ? _GEN_6452 : _GEN_6451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6454 = io_inputBit | _GEN_6453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6455 = i == 10'h183 ? _GEN_6454 : _GEN_6453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6456 = ~io_inputBit ? 1'h0 : _GEN_6455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6457 = i == 10'h184 ? _GEN_6456 : _GEN_6455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6458 = io_inputBit | _GEN_6457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6459 = i == 10'h184 ? _GEN_6458 : _GEN_6457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6460 = ~io_inputBit ? 1'h0 : _GEN_6459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6461 = i == 10'h185 ? _GEN_6460 : _GEN_6459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6462 = io_inputBit | _GEN_6461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6463 = i == 10'h185 ? _GEN_6462 : _GEN_6461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6464 = ~io_inputBit ? 1'h0 : _GEN_6463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6465 = i == 10'h186 ? _GEN_6464 : _GEN_6463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6466 = io_inputBit | _GEN_6465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6467 = i == 10'h186 ? _GEN_6466 : _GEN_6465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6468 = ~io_inputBit ? 1'h0 : _GEN_6467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6469 = i == 10'h187 ? _GEN_6468 : _GEN_6467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6470 = io_inputBit | _GEN_6469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6471 = i == 10'h187 ? _GEN_6470 : _GEN_6469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6472 = ~io_inputBit ? 1'h0 : _GEN_6471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6473 = i == 10'h188 ? _GEN_6472 : _GEN_6471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6474 = io_inputBit | _GEN_6473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6475 = i == 10'h188 ? _GEN_6474 : _GEN_6473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6476 = ~io_inputBit ? 1'h0 : _GEN_6475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6477 = i == 10'h189 ? _GEN_6476 : _GEN_6475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6478 = io_inputBit | _GEN_6477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6479 = i == 10'h189 ? _GEN_6478 : _GEN_6477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6480 = ~io_inputBit ? 1'h0 : _GEN_6479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6481 = i == 10'h18a ? _GEN_6480 : _GEN_6479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6482 = io_inputBit | _GEN_6481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6483 = i == 10'h18a ? _GEN_6482 : _GEN_6481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6484 = ~io_inputBit ? 1'h0 : _GEN_6483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6485 = i == 10'h18b ? _GEN_6484 : _GEN_6483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6486 = io_inputBit | _GEN_6485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6487 = i == 10'h18b ? _GEN_6486 : _GEN_6485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6488 = ~io_inputBit ? 1'h0 : _GEN_6487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6489 = i == 10'h18c ? _GEN_6488 : _GEN_6487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6490 = io_inputBit | _GEN_6489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6491 = i == 10'h18c ? _GEN_6490 : _GEN_6489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6492 = ~io_inputBit ? 1'h0 : _GEN_6491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6493 = i == 10'h18d ? _GEN_6492 : _GEN_6491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6494 = io_inputBit | _GEN_6493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6495 = i == 10'h18d ? _GEN_6494 : _GEN_6493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6496 = ~io_inputBit ? 1'h0 : _GEN_6495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6497 = i == 10'h18e ? _GEN_6496 : _GEN_6495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6498 = io_inputBit | _GEN_6497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6499 = i == 10'h18e ? _GEN_6498 : _GEN_6497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6500 = ~io_inputBit ? 1'h0 : _GEN_6499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6501 = i == 10'h18f ? _GEN_6500 : _GEN_6499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6502 = io_inputBit | _GEN_6501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6503 = i == 10'h18f ? _GEN_6502 : _GEN_6501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6504 = ~io_inputBit ? 1'h0 : _GEN_6503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6505 = i == 10'h190 ? _GEN_6504 : _GEN_6503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6506 = io_inputBit | _GEN_6505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6507 = i == 10'h190 ? _GEN_6506 : _GEN_6505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6508 = ~io_inputBit ? 1'h0 : _GEN_6507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6509 = i == 10'h191 ? _GEN_6508 : _GEN_6507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6510 = io_inputBit | _GEN_6509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6511 = i == 10'h191 ? _GEN_6510 : _GEN_6509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6512 = ~io_inputBit ? 1'h0 : _GEN_6511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6513 = i == 10'h192 ? _GEN_6512 : _GEN_6511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6514 = io_inputBit | _GEN_6513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6515 = i == 10'h192 ? _GEN_6514 : _GEN_6513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6516 = ~io_inputBit ? 1'h0 : _GEN_6515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6517 = i == 10'h193 ? _GEN_6516 : _GEN_6515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6518 = io_inputBit | _GEN_6517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6519 = i == 10'h193 ? _GEN_6518 : _GEN_6517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6520 = ~io_inputBit ? 1'h0 : _GEN_6519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6521 = i == 10'h194 ? _GEN_6520 : _GEN_6519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6522 = io_inputBit | _GEN_6521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6524 = ~io_inputBit ? 1'h0 : _GEN_6173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6525 = i == 10'h1 ? _GEN_6524 : _GEN_6173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6526 = io_inputBit ? 1'h0 : _GEN_6525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6527 = i == 10'h2 ? _GEN_6526 : _GEN_6525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6528 = ~io_inputBit ? 1'h0 : _GEN_6527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6529 = i == 10'h4 ? _GEN_6528 : _GEN_6527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6530 = io_inputBit ? 1'h0 : _GEN_6529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6531 = i == 10'h5 ? _GEN_6530 : _GEN_6529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6532 = ~io_inputBit ? 1'h0 : _GEN_6531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6533 = i == 10'ha ? _GEN_6532 : _GEN_6531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6534 = ~io_inputBit ? 1'h0 : _GEN_6533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6535 = i == 10'h16 ? _GEN_6534 : _GEN_6533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6536 = io_inputBit ? 1'h0 : _GEN_6535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6537 = i == 10'h18 ? _GEN_6536 : _GEN_6535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6538 = ~io_inputBit ? 1'h0 : _GEN_6537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6539 = i == 10'h2e ? _GEN_6538 : _GEN_6537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6540 = io_inputBit ? 1'h0 : _GEN_6539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6541 = i == 10'h64 ? _GEN_6540 : _GEN_6539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6542 = ~io_inputBit ? 1'h0 : _GEN_6541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6543 = i == 10'hbd ? _GEN_6542 : _GEN_6541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6544 = ~io_inputBit ? 1'h0 : _GEN_6543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6545 = i == 10'h2f9 ? _GEN_6544 : _GEN_6543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6546 = io_inputBit | _GEN_6545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6547 = i == 10'h2f9 ? _GEN_6546 : _GEN_6545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6548 = ~io_inputBit ? 1'h0 : _GEN_6547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6549 = i == 10'h2fa ? _GEN_6548 : _GEN_6547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6550 = io_inputBit | _GEN_6549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6551 = i == 10'h2fa ? _GEN_6550 : _GEN_6549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6552 = ~io_inputBit ? 1'h0 : _GEN_6551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6553 = i == 10'h2fb ? _GEN_6552 : _GEN_6551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6554 = io_inputBit | _GEN_6553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6555 = i == 10'h2fb ? _GEN_6554 : _GEN_6553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6556 = ~io_inputBit ? 1'h0 : _GEN_6555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6557 = i == 10'h2fc ? _GEN_6556 : _GEN_6555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6558 = io_inputBit | _GEN_6557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6559 = i == 10'h2fc ? _GEN_6558 : _GEN_6557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6560 = ~io_inputBit ? 1'h0 : _GEN_6559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6561 = i == 10'h2fd ? _GEN_6560 : _GEN_6559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6562 = io_inputBit | _GEN_6561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6563 = i == 10'h2fd ? _GEN_6562 : _GEN_6561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6564 = ~io_inputBit ? 1'h0 : _GEN_6563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6565 = i == 10'h2fe ? _GEN_6564 : _GEN_6563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6566 = io_inputBit | _GEN_6565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6567 = i == 10'h2fe ? _GEN_6566 : _GEN_6565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6568 = ~io_inputBit ? 1'h0 : _GEN_6567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6569 = i == 10'h2ff ? _GEN_6568 : _GEN_6567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6570 = io_inputBit | _GEN_6569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6571 = i == 10'h2ff ? _GEN_6570 : _GEN_6569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6572 = ~io_inputBit ? 1'h0 : _GEN_6571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6573 = i == 10'h300 ? _GEN_6572 : _GEN_6571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6574 = io_inputBit | _GEN_6573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6575 = i == 10'h300 ? _GEN_6574 : _GEN_6573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6576 = ~io_inputBit ? 1'h0 : _GEN_6575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6577 = i == 10'h301 ? _GEN_6576 : _GEN_6575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6578 = io_inputBit | _GEN_6577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6579 = i == 10'h301 ? _GEN_6578 : _GEN_6577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6580 = ~io_inputBit ? 1'h0 : _GEN_6579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6581 = i == 10'h302 ? _GEN_6580 : _GEN_6579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6582 = io_inputBit | _GEN_6581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6583 = i == 10'h302 ? _GEN_6582 : _GEN_6581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6584 = ~io_inputBit ? 1'h0 : _GEN_6583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6585 = i == 10'h303 ? _GEN_6584 : _GEN_6583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6586 = io_inputBit | _GEN_6585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6587 = i == 10'h303 ? _GEN_6586 : _GEN_6585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6588 = ~io_inputBit ? 1'h0 : _GEN_6587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6589 = i == 10'h304 ? _GEN_6588 : _GEN_6587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6590 = io_inputBit | _GEN_6589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6591 = i == 10'h304 ? _GEN_6590 : _GEN_6589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6592 = ~io_inputBit ? 1'h0 : _GEN_6591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6593 = i == 10'h305 ? _GEN_6592 : _GEN_6591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6594 = io_inputBit | _GEN_6593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6595 = i == 10'h305 ? _GEN_6594 : _GEN_6593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6596 = ~io_inputBit ? 1'h0 : _GEN_6595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6597 = i == 10'h306 ? _GEN_6596 : _GEN_6595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6598 = io_inputBit | _GEN_6597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6599 = i == 10'h306 ? _GEN_6598 : _GEN_6597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6600 = ~io_inputBit ? 1'h0 : _GEN_6599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6601 = i == 10'h307 ? _GEN_6600 : _GEN_6599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6602 = io_inputBit | _GEN_6601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6603 = i == 10'h307 ? _GEN_6602 : _GEN_6601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6604 = ~io_inputBit ? 1'h0 : _GEN_6603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6605 = i == 10'h308 ? _GEN_6604 : _GEN_6603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6606 = io_inputBit | _GEN_6605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6607 = i == 10'h308 ? _GEN_6606 : _GEN_6605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6608 = ~io_inputBit ? 1'h0 : _GEN_6607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6609 = i == 10'h309 ? _GEN_6608 : _GEN_6607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6610 = io_inputBit | _GEN_6609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6611 = i == 10'h309 ? _GEN_6610 : _GEN_6609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6612 = ~io_inputBit ? 1'h0 : _GEN_6611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6613 = i == 10'h30a ? _GEN_6612 : _GEN_6611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6614 = io_inputBit | _GEN_6613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6615 = i == 10'h30a ? _GEN_6614 : _GEN_6613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6616 = ~io_inputBit ? 1'h0 : _GEN_6615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6617 = i == 10'h30b ? _GEN_6616 : _GEN_6615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6618 = io_inputBit | _GEN_6617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6619 = i == 10'h30b ? _GEN_6618 : _GEN_6617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6620 = ~io_inputBit ? 1'h0 : _GEN_6619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6621 = i == 10'h30c ? _GEN_6620 : _GEN_6619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6622 = io_inputBit | _GEN_6621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6623 = i == 10'h30c ? _GEN_6622 : _GEN_6621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6624 = ~io_inputBit ? 1'h0 : _GEN_6623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6625 = i == 10'h30d ? _GEN_6624 : _GEN_6623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6626 = io_inputBit | _GEN_6625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6627 = i == 10'h30d ? _GEN_6626 : _GEN_6625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6628 = ~io_inputBit ? 1'h0 : _GEN_6627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6629 = i == 10'h30e ? _GEN_6628 : _GEN_6627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6630 = io_inputBit | _GEN_6629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6631 = i == 10'h30e ? _GEN_6630 : _GEN_6629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6632 = ~io_inputBit ? 1'h0 : _GEN_6631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6633 = i == 10'h30f ? _GEN_6632 : _GEN_6631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6634 = io_inputBit | _GEN_6633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6635 = i == 10'h30f ? _GEN_6634 : _GEN_6633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6636 = ~io_inputBit ? 1'h0 : _GEN_6635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6637 = i == 10'h310 ? _GEN_6636 : _GEN_6635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6638 = io_inputBit | _GEN_6637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6639 = i == 10'h310 ? _GEN_6638 : _GEN_6637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6640 = ~io_inputBit ? 1'h0 : _GEN_6639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6641 = i == 10'h311 ? _GEN_6640 : _GEN_6639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6642 = io_inputBit | _GEN_6641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6643 = i == 10'h311 ? _GEN_6642 : _GEN_6641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6644 = ~io_inputBit ? 1'h0 : _GEN_6643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6645 = i == 10'h312 ? _GEN_6644 : _GEN_6643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6646 = io_inputBit | _GEN_6645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6647 = i == 10'h312 ? _GEN_6646 : _GEN_6645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6648 = ~io_inputBit ? 1'h0 : _GEN_6647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6649 = i == 10'h313 ? _GEN_6648 : _GEN_6647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6650 = io_inputBit | _GEN_6649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6651 = i == 10'h313 ? _GEN_6650 : _GEN_6649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6652 = ~io_inputBit ? 1'h0 : _GEN_6651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6653 = i == 10'h314 ? _GEN_6652 : _GEN_6651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6654 = io_inputBit | _GEN_6653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6655 = i == 10'h314 ? _GEN_6654 : _GEN_6653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6656 = ~io_inputBit ? 1'h0 : _GEN_6655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6657 = i == 10'h315 ? _GEN_6656 : _GEN_6655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6658 = io_inputBit | _GEN_6657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6659 = i == 10'h315 ? _GEN_6658 : _GEN_6657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6660 = ~io_inputBit ? 1'h0 : _GEN_6659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6661 = i == 10'h316 ? _GEN_6660 : _GEN_6659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6662 = io_inputBit | _GEN_6661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6663 = i == 10'h316 ? _GEN_6662 : _GEN_6661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6664 = ~io_inputBit ? 1'h0 : _GEN_6663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6665 = i == 10'h317 ? _GEN_6664 : _GEN_6663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6666 = io_inputBit | _GEN_6665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6667 = i == 10'h317 ? _GEN_6666 : _GEN_6665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6668 = ~io_inputBit ? 1'h0 : _GEN_6667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6669 = i == 10'h318 ? _GEN_6668 : _GEN_6667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6670 = io_inputBit | _GEN_6669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6671 = i == 10'h318 ? _GEN_6670 : _GEN_6669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6672 = ~io_inputBit ? 1'h0 : _GEN_6671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6673 = i == 10'h319 ? _GEN_6672 : _GEN_6671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6674 = io_inputBit | _GEN_6673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6675 = i == 10'h319 ? _GEN_6674 : _GEN_6673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6676 = ~io_inputBit ? 1'h0 : _GEN_6675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6677 = i == 10'h31a ? _GEN_6676 : _GEN_6675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6678 = io_inputBit | _GEN_6677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6679 = i == 10'h31a ? _GEN_6678 : _GEN_6677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6680 = ~io_inputBit ? 1'h0 : _GEN_6679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6681 = i == 10'h31b ? _GEN_6680 : _GEN_6679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6682 = io_inputBit | _GEN_6681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6683 = i == 10'h31b ? _GEN_6682 : _GEN_6681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6684 = ~io_inputBit ? 1'h0 : _GEN_6683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6685 = i == 10'h31c ? _GEN_6684 : _GEN_6683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6686 = io_inputBit | _GEN_6685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6687 = i == 10'h31c ? _GEN_6686 : _GEN_6685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6688 = ~io_inputBit ? 1'h0 : _GEN_6687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6689 = i == 10'h31d ? _GEN_6688 : _GEN_6687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6690 = io_inputBit | _GEN_6689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6691 = i == 10'h31d ? _GEN_6690 : _GEN_6689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6692 = ~io_inputBit ? 1'h0 : _GEN_6691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6693 = i == 10'h31e ? _GEN_6692 : _GEN_6691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6694 = io_inputBit | _GEN_6693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6695 = i == 10'h31e ? _GEN_6694 : _GEN_6693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6696 = ~io_inputBit ? 1'h0 : _GEN_6695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6697 = i == 10'h31f ? _GEN_6696 : _GEN_6695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6698 = io_inputBit | _GEN_6697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6699 = i == 10'h31f ? _GEN_6698 : _GEN_6697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6700 = ~io_inputBit ? 1'h0 : _GEN_6699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6701 = i == 10'h320 ? _GEN_6700 : _GEN_6699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6702 = io_inputBit | _GEN_6701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6703 = i == 10'h320 ? _GEN_6702 : _GEN_6701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6704 = ~io_inputBit ? 1'h0 : _GEN_6703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6705 = i == 10'h321 ? _GEN_6704 : _GEN_6703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6706 = io_inputBit | _GEN_6705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6707 = i == 10'h321 ? _GEN_6706 : _GEN_6705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6708 = ~io_inputBit ? 1'h0 : _GEN_6707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6709 = i == 10'h322 ? _GEN_6708 : _GEN_6707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6710 = io_inputBit | _GEN_6709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6711 = i == 10'h322 ? _GEN_6710 : _GEN_6709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6712 = ~io_inputBit ? 1'h0 : _GEN_6711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6713 = i == 10'h323 ? _GEN_6712 : _GEN_6711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6714 = io_inputBit | _GEN_6713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6715 = i == 10'h323 ? _GEN_6714 : _GEN_6713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6716 = ~io_inputBit ? 1'h0 : _GEN_6715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6717 = i == 10'h324 ? _GEN_6716 : _GEN_6715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6718 = io_inputBit | _GEN_6717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6719 = i == 10'h324 ? _GEN_6718 : _GEN_6717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6720 = ~io_inputBit ? 1'h0 : _GEN_6719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6721 = i == 10'h325 ? _GEN_6720 : _GEN_6719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6722 = io_inputBit | _GEN_6721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6723 = i == 10'h325 ? _GEN_6722 : _GEN_6721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6724 = ~io_inputBit ? 1'h0 : _GEN_6723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6725 = i == 10'h326 ? _GEN_6724 : _GEN_6723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6726 = io_inputBit | _GEN_6725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6727 = i == 10'h326 ? _GEN_6726 : _GEN_6725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6728 = ~io_inputBit ? 1'h0 : _GEN_6727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6729 = i == 10'h327 ? _GEN_6728 : _GEN_6727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6730 = io_inputBit | _GEN_6729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6731 = i == 10'h327 ? _GEN_6730 : _GEN_6729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6732 = ~io_inputBit ? 1'h0 : _GEN_6731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6733 = i == 10'h328 ? _GEN_6732 : _GEN_6731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6734 = io_inputBit | _GEN_6733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6735 = i == 10'h328 ? _GEN_6734 : _GEN_6733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6736 = ~io_inputBit ? 1'h0 : _GEN_6735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6737 = i == 10'h329 ? _GEN_6736 : _GEN_6735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6738 = io_inputBit | _GEN_6737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6739 = i == 10'h329 ? _GEN_6738 : _GEN_6737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6740 = ~io_inputBit ? 1'h0 : _GEN_6739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_6741 = i == 10'h32a ? _GEN_6740 : _GEN_6739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_6742 = io_inputBit | _GEN_6741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _T_6747 = counter < 5'h11; // @[lut_mem_online.scala 248:22]
  wire  _T_6749 = counter >= 5'ha; // @[lut_mem_online.scala 256:30]
  wire [4:0] _outResult_T_1 = counter - 5'ha; // @[lut_mem_online.scala 258:41]
  wire  _GEN_6752 = 4'h1 == _outResult_T_1[3:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6753 = 4'h2 == _outResult_T_1[3:0] ? buffer_2 : _GEN_6752; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6754 = 4'h3 == _outResult_T_1[3:0] ? buffer_3 : _GEN_6753; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6755 = 4'h4 == _outResult_T_1[3:0] ? buffer_4 : _GEN_6754; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6756 = 4'h5 == _outResult_T_1[3:0] ? buffer_5 : _GEN_6755; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6757 = 4'h6 == _outResult_T_1[3:0] ? buffer_6 : _GEN_6756; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6758 = 4'h7 == _outResult_T_1[3:0] ? 1'h0 : _GEN_6757; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6759 = 4'h8 == _outResult_T_1[3:0] ? 1'h0 : _GEN_6758; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_6760 = 4'h9 == _outResult_T_1[3:0] ? 1'h0 : _GEN_6759; // @[lut_mem_online.scala 258:{23,23}]
  wire  _T_6753 = ~reset; // @[lut_mem_online.scala 260:21]
  wire  _GEN_6762 = counter >= 5'ha ? _GEN_6760 : outResult; // @[lut_mem_online.scala 256:42 258:23 214:26]
  wire  _GEN_6764 = _T_2 ? 1'h0 : _GEN_6762; // @[lut_mem_online.scala 253:35 255:23]
  wire  _T_6754 = i < 10'h1ff; // @[lut_mem_online.scala 271:18]
  wire [11:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 281:24]
  wire [11:0] _i_T_2 = _i_T + 12'h1; // @[lut_mem_online.scala 281:28]
  wire [11:0] _i_T_5 = _i_T + 12'h2; // @[lut_mem_online.scala 283:28]
  wire [11:0] _GEN_6765 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 282:45 283:17 205:18]
  wire [11:0] _GEN_6766 = _T_10 ? _i_T_2 : _GEN_6765; // @[lut_mem_online.scala 280:39 281:17]
  wire  _T_6759 = i < 10'h3ff; // @[lut_mem_online.scala 286:24]
  wire [9:0] _GEN_6767 = i < 10'h3ff ? 10'h3ff : i; // @[lut_mem_online.scala 286:63 294:15 205:18]
  wire [11:0] _GEN_6768 = i < 10'h1ff ? _GEN_6766 : {{2'd0}, _GEN_6767}; // @[lut_mem_online.scala 271:61]
  wire [4:0] _counter_T_1 = counter + 5'h1; // @[lut_mem_online.scala 297:30]
  wire  _GEN_6770 = counter < 5'h11 & _GEN_6764; // @[lut_mem_online.scala 248:52 300:21]
  wire [11:0] _GEN_6771 = counter < 5'h11 ? _GEN_6768 : {{2'd0}, i}; // @[lut_mem_online.scala 205:18 248:52]
  wire  _GEN_6794 = io_start & _GEN_6770; // @[lut_mem_online.scala 219:29 323:15]
  wire [11:0] _GEN_6795 = io_start ? _GEN_6771 : 12'h0; // @[lut_mem_online.scala 219:29 321:7]
  wire [11:0] _GEN_6798 = reset ? 12'h0 : _GEN_6795; // @[lut_mem_online.scala 205:{18,18}]
  wire  _GEN_6799 = io_start & _T_6747; // @[lut_mem_online.scala 260:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 330:16]
  always @(posedge clock) begin
    i <= _GEN_6798[9:0]; // @[lut_mem_online.scala 205:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'hc5) begin // @[lut_mem_online.scala 234:34]
          buffer_0 <= _GEN_6190;
        end else if (i == 10'hc5) begin // @[lut_mem_online.scala 234:34]
          buffer_0 <= _GEN_6188;
        end else begin
          buffer_0 <= _GEN_6187;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 234:34]
          buffer_1 <= _GEN_6222;
        end else if (i == 10'hc9) begin // @[lut_mem_online.scala 234:34]
          buffer_1 <= _GEN_6220;
        end else begin
          buffer_1 <= _GEN_6219;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_2 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_2 <= _GEN_6265;
          end
        end else begin
          buffer_2 <= _GEN_6265;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_3 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_3 <= _GEN_6333;
          end
        end else begin
          buffer_3 <= _GEN_6333;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'hc9) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_4 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_4 <= _GEN_6401;
          end
        end else begin
          buffer_4 <= _GEN_6401;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'h194) begin // @[lut_mem_online.scala 234:34]
          buffer_5 <= _GEN_6522;
        end else if (i == 10'h194) begin // @[lut_mem_online.scala 234:34]
          buffer_5 <= _GEN_6520;
        end else begin
          buffer_5 <= _GEN_6519;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'ha) begin // @[lut_mem_online.scala 231:36]
        if (i == 10'h32a) begin // @[lut_mem_online.scala 234:34]
          buffer_6 <= _GEN_6742;
        end else if (i == 10'h32a) begin // @[lut_mem_online.scala 234:34]
          buffer_6 <= _GEN_6740;
        end else begin
          buffer_6 <= _GEN_6739;
        end
      end
    end
    if (reset) begin // @[lut_mem_online.scala 211:24]
      counter <= 5'h0; // @[lut_mem_online.scala 211:24]
    end else if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 5'h11) begin // @[lut_mem_online.scala 248:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 297:19]
      end
    end else begin
      counter <= 5'h0; // @[lut_mem_online.scala 322:13]
    end
    if (reset) begin // @[lut_mem_online.scala 214:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 214:26]
    end else begin
      outResult <= _GEN_6794;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_6747 & ~_T_2 & _T_6749 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 260:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_6799 & _T_6754 & _T_6753) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 274:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_6799 & ~_T_6754 & _T_6759 & _T_6753) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 289:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
