module LutMembershipFunctionOnline_8(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [7:0] i; // @[lut_mem_online.scala 206:18]
  reg  buffer_0; // @[lut_mem_online.scala 210:19]
  reg  buffer_1; // @[lut_mem_online.scala 210:19]
  reg  buffer_2; // @[lut_mem_online.scala 210:19]
  reg  buffer_3; // @[lut_mem_online.scala 210:19]
  reg  buffer_4; // @[lut_mem_online.scala 210:19]
  reg  buffer_5; // @[lut_mem_online.scala 210:19]
  reg  buffer_6; // @[lut_mem_online.scala 210:19]
  reg [4:0] counter; // @[lut_mem_online.scala 212:24]
  reg  outResult; // @[lut_mem_online.scala 215:26]
  wire  _GEN_0 = i == 8'h0 ? 1'h0 : buffer_0; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_1 = i == 8'h1 ? 1'h0 : _GEN_0; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2 = i == 8'h3 ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_4 = i == 8'h10 ? 1'h0 : i == 8'h7 | _GEN_2; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_6 = i == 8'h44 ? 1'h0 : i == 8'h21 | _GEN_4; // @[lut_mem_online.scala 235:34 239:30]
  wire [8:0] _GEN_3306 = {{1'd0}, i}; // @[lut_mem_online.scala 235:20]
  wire [9:0] _GEN_3307 = {{2'd0}, i}; // @[lut_mem_online.scala 235:20]
  wire  _GEN_10 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_3307 == 10'h22a | (_GEN_3306 == 9'h114 | (i == 8'h89 | _GEN_6)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_11 = i == 8'h0 ? 1'h0 : buffer_1; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_12 = i == 8'h1 ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_13 = i == 8'h3 ? 1'h0 : _GEN_12; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_16 = i == 8'h21 ? 1'h0 : i == 8'h20 | (i == 8'hf | _GEN_13); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_18 = i == 8'h42 ? 1'h0 : i == 8'h22 | _GEN_16; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_20 = i == 8'h46 ? 1'h0 : i == 8'h44 | _GEN_18; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_22 = i == 8'h89 ? 1'h0 : i == 8'h85 | _GEN_20; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_25 = _GEN_3306 == 9'h114 ? 1'h0 : _GEN_3306 == 9'h10c | (i == 8'h8d | _GEN_22); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_28 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_3307 == 10'h21a | (_GEN_3306 == 9'h11c | _GEN_25); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_29 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_28; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_32 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_3307 == 10'h23a | (_GEN_3307 == 10'h22a | _GEN_29); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_33 = i == 8'h0 ? 1'h0 : buffer_2; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_34 = i == 8'h1 ? 1'h0 : _GEN_33; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_35 = i == 8'h8 ? 1'h0 : _GEN_34; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_36 = i == 8'hf ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_37 = i == 8'h11 ? 1'h0 : _GEN_36; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_38 = i == 8'h20 ? 1'h0 : _GEN_37; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_39 = i == 8'h23 ? 1'h0 : _GEN_38; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_41 = i == 8'h43 ? 1'h0 : i == 8'h42 | _GEN_39; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_43 = i == 8'h45 ? 1'h0 : i == 8'h44 | _GEN_41; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_45 = i == 8'h47 ? 1'h0 : i == 8'h46 | _GEN_43; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_46 = i == 8'h85 ? 1'h0 : _GEN_45; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_48 = i == 8'h89 ? 1'h0 : i == 8'h87 | _GEN_46; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_50 = i == 8'h8d ? 1'h0 : i == 8'h8b | _GEN_48; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_52 = _GEN_3306 == 9'h10c ? 1'h0 : i == 8'h8f | _GEN_50; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_54 = _GEN_3306 == 9'h114 ? 1'h0 : _GEN_3306 == 9'h110 | _GEN_52; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_56 = _GEN_3306 == 9'h11c ? 1'h0 : _GEN_3306 == 9'h118 | _GEN_54; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_58 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_3306 == 9'h120 | _GEN_56; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_61 = _GEN_3307 == 10'h222 ? 1'h0 : _GEN_3307 == 10'h222 | (_GEN_3307 == 10'h21a | _GEN_58); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_62 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_61; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_65 = _GEN_3307 == 10'h232 ? 1'h0 : _GEN_3307 == 10'h232 | (_GEN_3307 == 10'h22a | _GEN_62); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_66 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_65; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_69 = _GEN_3307 == 10'h242 ? 1'h0 : _GEN_3307 == 10'h242 | (_GEN_3307 == 10'h23a | _GEN_66); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_70 = i == 8'h0 ? 1'h0 : buffer_3; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_71 = i == 8'h1 ? 1'h0 : _GEN_70; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_72 = i == 8'h8 ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_73 = i == 8'hf ? 1'h0 : _GEN_72; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_74 = i == 8'h11 ? 1'h0 : _GEN_73; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_75 = i == 8'h20 ? 1'h0 : _GEN_74; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_76 = i == 8'h23 ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_77 = i == 8'h85 ? 1'h0 : _GEN_76; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_79 = i == 8'h87 ? 1'h0 : i == 8'h86 | _GEN_77; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_81 = i == 8'h89 ? 1'h0 : i == 8'h88 | _GEN_79; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_83 = i == 8'h8b ? 1'h0 : i == 8'h8a | _GEN_81; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_85 = i == 8'h8d ? 1'h0 : i == 8'h8c | _GEN_83; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_87 = i == 8'h8f ? 1'h0 : i == 8'h8e | _GEN_85; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_89 = _GEN_3306 == 9'h10c ? 1'h0 : i == 8'h90 | _GEN_87; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_91 = _GEN_3306 == 9'h110 ? 1'h0 : _GEN_3306 == 9'h10e | _GEN_89; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_93 = _GEN_3306 == 9'h114 ? 1'h0 : _GEN_3306 == 9'h112 | _GEN_91; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_95 = _GEN_3306 == 9'h118 ? 1'h0 : _GEN_3306 == 9'h116 | _GEN_93; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_97 = _GEN_3306 == 9'h11c ? 1'h0 : _GEN_3306 == 9'h11a | _GEN_95; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_99 = _GEN_3306 == 9'h120 ? 1'h0 : _GEN_3306 == 9'h11e | _GEN_97; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_101 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_3306 == 9'h122 | _GEN_99; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_104 = _GEN_3307 == 10'h21e ? 1'h0 : _GEN_3307 == 10'h21e | (_GEN_3307 == 10'h21a | _GEN_101); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_105 = _GEN_3307 == 10'h222 ? 1'h0 : _GEN_104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_108 = _GEN_3307 == 10'h226 ? 1'h0 : _GEN_3307 == 10'h226 | (_GEN_3307 == 10'h222 | _GEN_105); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_109 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_108; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_112 = _GEN_3307 == 10'h22e ? 1'h0 : _GEN_3307 == 10'h22e | (_GEN_3307 == 10'h22a | _GEN_109); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_113 = _GEN_3307 == 10'h232 ? 1'h0 : _GEN_112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_116 = _GEN_3307 == 10'h236 ? 1'h0 : _GEN_3307 == 10'h236 | (_GEN_3307 == 10'h232 | _GEN_113); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_117 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_120 = _GEN_3307 == 10'h23e ? 1'h0 : _GEN_3307 == 10'h23e | (_GEN_3307 == 10'h23a | _GEN_117); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_121 = _GEN_3307 == 10'h242 ? 1'h0 : _GEN_120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_124 = _GEN_3307 == 10'h246 ? 1'h0 : _GEN_3307 == 10'h246 | (_GEN_3307 == 10'h242 | _GEN_121); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_125 = i == 8'h0 ? 1'h0 : buffer_4; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_126 = i == 8'h1 ? 1'h0 : _GEN_125; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_127 = i == 8'h8 ? 1'h0 : _GEN_126; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_129 = i == 8'h11 ? 1'h0 : i == 8'hf | _GEN_127; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_131 = i == 8'h48 ? 1'h0 : i == 8'h20 | _GEN_129; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_132 = i == 8'h91 ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_134 = _GEN_3306 == 9'h10c ? 1'h0 : _GEN_3306 == 9'h10b | _GEN_132; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_136 = _GEN_3306 == 9'h10e ? 1'h0 : _GEN_3306 == 9'h10d | _GEN_134; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_138 = _GEN_3306 == 9'h110 ? 1'h0 : _GEN_3306 == 9'h10f | _GEN_136; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_140 = _GEN_3306 == 9'h112 ? 1'h0 : _GEN_3306 == 9'h111 | _GEN_138; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_142 = _GEN_3306 == 9'h114 ? 1'h0 : _GEN_3306 == 9'h113 | _GEN_140; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_144 = _GEN_3306 == 9'h116 ? 1'h0 : _GEN_3306 == 9'h115 | _GEN_142; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_146 = _GEN_3306 == 9'h118 ? 1'h0 : _GEN_3306 == 9'h117 | _GEN_144; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_148 = _GEN_3306 == 9'h11a ? 1'h0 : _GEN_3306 == 9'h119 | _GEN_146; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_150 = _GEN_3306 == 9'h11c ? 1'h0 : _GEN_3306 == 9'h11b | _GEN_148; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_152 = _GEN_3306 == 9'h11e ? 1'h0 : _GEN_3306 == 9'h11d | _GEN_150; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_154 = _GEN_3306 == 9'h120 ? 1'h0 : _GEN_3306 == 9'h11f | _GEN_152; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_156 = _GEN_3306 == 9'h122 ? 1'h0 : _GEN_3306 == 9'h121 | _GEN_154; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_159 = _GEN_3307 == 10'h218 ? 1'h0 : _GEN_3307 == 10'h218 | (_GEN_3306 == 9'h123 | _GEN_156); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_160 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_159; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_163 = _GEN_3307 == 10'h21c ? 1'h0 : _GEN_3307 == 10'h21c | (_GEN_3307 == 10'h21a | _GEN_160); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_164 = _GEN_3307 == 10'h21e ? 1'h0 : _GEN_163; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_167 = _GEN_3307 == 10'h220 ? 1'h0 : _GEN_3307 == 10'h220 | (_GEN_3307 == 10'h21e | _GEN_164); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_168 = _GEN_3307 == 10'h222 ? 1'h0 : _GEN_167; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_171 = _GEN_3307 == 10'h224 ? 1'h0 : _GEN_3307 == 10'h224 | (_GEN_3307 == 10'h222 | _GEN_168); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_172 = _GEN_3307 == 10'h226 ? 1'h0 : _GEN_171; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_175 = _GEN_3307 == 10'h228 ? 1'h0 : _GEN_3307 == 10'h228 | (_GEN_3307 == 10'h226 | _GEN_172); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_176 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_175; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_179 = _GEN_3307 == 10'h22c ? 1'h0 : _GEN_3307 == 10'h22c | (_GEN_3307 == 10'h22a | _GEN_176); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_180 = _GEN_3307 == 10'h22e ? 1'h0 : _GEN_179; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_183 = _GEN_3307 == 10'h230 ? 1'h0 : _GEN_3307 == 10'h230 | (_GEN_3307 == 10'h22e | _GEN_180); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_184 = _GEN_3307 == 10'h232 ? 1'h0 : _GEN_183; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_187 = _GEN_3307 == 10'h234 ? 1'h0 : _GEN_3307 == 10'h234 | (_GEN_3307 == 10'h232 | _GEN_184); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_188 = _GEN_3307 == 10'h236 ? 1'h0 : _GEN_187; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_191 = _GEN_3307 == 10'h238 ? 1'h0 : _GEN_3307 == 10'h238 | (_GEN_3307 == 10'h236 | _GEN_188); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_192 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_191; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_195 = _GEN_3307 == 10'h23c ? 1'h0 : _GEN_3307 == 10'h23c | (_GEN_3307 == 10'h23a | _GEN_192); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_196 = _GEN_3307 == 10'h23e ? 1'h0 : _GEN_195; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_199 = _GEN_3307 == 10'h240 ? 1'h0 : _GEN_3307 == 10'h240 | (_GEN_3307 == 10'h23e | _GEN_196); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_200 = _GEN_3307 == 10'h242 ? 1'h0 : _GEN_199; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_203 = _GEN_3307 == 10'h244 ? 1'h0 : _GEN_3307 == 10'h244 | (_GEN_3307 == 10'h242 | _GEN_200); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_204 = _GEN_3307 == 10'h246 ? 1'h0 : _GEN_203; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_207 = _GEN_3307 == 10'h248 ? 1'h0 : _GEN_3307 == 10'h248 | (_GEN_3307 == 10'h246 | _GEN_204); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_208 = i == 8'h0 ? 1'h0 : buffer_5; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_209 = i == 8'h1 ? 1'h0 : _GEN_208; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_210 = i == 8'h8 ? 1'h0 : _GEN_209; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_211 = i == 8'hf ? 1'h0 : _GEN_210; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_212 = i == 8'h11 ? 1'h0 : _GEN_211; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_213 = i == 8'h20 ? 1'h0 : _GEN_212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_214 = i == 8'h48 ? 1'h0 : _GEN_213; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_215 = _GEN_3306 == 9'h10b ? 1'h0 : _GEN_214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_216 = _GEN_3306 == 9'h124 ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_217 = _GEN_3307 == 10'h218 ? 1'h0 : _GEN_216; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_220 = _GEN_3307 == 10'h219 ? 1'h0 : _GEN_3307 == 10'h219 | (_GEN_3307 == 10'h218 | _GEN_217); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_221 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_224 = _GEN_3307 == 10'h21b ? 1'h0 : _GEN_3307 == 10'h21b | (_GEN_3307 == 10'h21a | _GEN_221); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_225 = _GEN_3307 == 10'h21c ? 1'h0 : _GEN_224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_228 = _GEN_3307 == 10'h21d ? 1'h0 : _GEN_3307 == 10'h21d | (_GEN_3307 == 10'h21c | _GEN_225); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_229 = _GEN_3307 == 10'h21e ? 1'h0 : _GEN_228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_232 = _GEN_3307 == 10'h21f ? 1'h0 : _GEN_3307 == 10'h21f | (_GEN_3307 == 10'h21e | _GEN_229); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_233 = _GEN_3307 == 10'h220 ? 1'h0 : _GEN_232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_236 = _GEN_3307 == 10'h221 ? 1'h0 : _GEN_3307 == 10'h221 | (_GEN_3307 == 10'h220 | _GEN_233); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_237 = _GEN_3307 == 10'h222 ? 1'h0 : _GEN_236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_240 = _GEN_3307 == 10'h223 ? 1'h0 : _GEN_3307 == 10'h223 | (_GEN_3307 == 10'h222 | _GEN_237); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_241 = _GEN_3307 == 10'h224 ? 1'h0 : _GEN_240; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_244 = _GEN_3307 == 10'h225 ? 1'h0 : _GEN_3307 == 10'h225 | (_GEN_3307 == 10'h224 | _GEN_241); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_245 = _GEN_3307 == 10'h226 ? 1'h0 : _GEN_244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_248 = _GEN_3307 == 10'h227 ? 1'h0 : _GEN_3307 == 10'h227 | (_GEN_3307 == 10'h226 | _GEN_245); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_249 = _GEN_3307 == 10'h228 ? 1'h0 : _GEN_248; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_252 = _GEN_3307 == 10'h229 ? 1'h0 : _GEN_3307 == 10'h229 | (_GEN_3307 == 10'h228 | _GEN_249); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_253 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_252; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_256 = _GEN_3307 == 10'h22b ? 1'h0 : _GEN_3307 == 10'h22b | (_GEN_3307 == 10'h22a | _GEN_253); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_257 = _GEN_3307 == 10'h22c ? 1'h0 : _GEN_256; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_260 = _GEN_3307 == 10'h22d ? 1'h0 : _GEN_3307 == 10'h22d | (_GEN_3307 == 10'h22c | _GEN_257); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_261 = _GEN_3307 == 10'h22e ? 1'h0 : _GEN_260; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_264 = _GEN_3307 == 10'h22f ? 1'h0 : _GEN_3307 == 10'h22f | (_GEN_3307 == 10'h22e | _GEN_261); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_265 = _GEN_3307 == 10'h230 ? 1'h0 : _GEN_264; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_268 = _GEN_3307 == 10'h231 ? 1'h0 : _GEN_3307 == 10'h231 | (_GEN_3307 == 10'h230 | _GEN_265); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_269 = _GEN_3307 == 10'h232 ? 1'h0 : _GEN_268; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_272 = _GEN_3307 == 10'h233 ? 1'h0 : _GEN_3307 == 10'h233 | (_GEN_3307 == 10'h232 | _GEN_269); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_273 = _GEN_3307 == 10'h234 ? 1'h0 : _GEN_272; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_276 = _GEN_3307 == 10'h235 ? 1'h0 : _GEN_3307 == 10'h235 | (_GEN_3307 == 10'h234 | _GEN_273); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_277 = _GEN_3307 == 10'h236 ? 1'h0 : _GEN_276; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_280 = _GEN_3307 == 10'h237 ? 1'h0 : _GEN_3307 == 10'h237 | (_GEN_3307 == 10'h236 | _GEN_277); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_281 = _GEN_3307 == 10'h238 ? 1'h0 : _GEN_280; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_284 = _GEN_3307 == 10'h239 ? 1'h0 : _GEN_3307 == 10'h239 | (_GEN_3307 == 10'h238 | _GEN_281); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_285 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_284; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_288 = _GEN_3307 == 10'h23b ? 1'h0 : _GEN_3307 == 10'h23b | (_GEN_3307 == 10'h23a | _GEN_285); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_289 = _GEN_3307 == 10'h23c ? 1'h0 : _GEN_288; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_292 = _GEN_3307 == 10'h23d ? 1'h0 : _GEN_3307 == 10'h23d | (_GEN_3307 == 10'h23c | _GEN_289); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_293 = _GEN_3307 == 10'h23e ? 1'h0 : _GEN_292; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_296 = _GEN_3307 == 10'h23f ? 1'h0 : _GEN_3307 == 10'h23f | (_GEN_3307 == 10'h23e | _GEN_293); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_297 = _GEN_3307 == 10'h240 ? 1'h0 : _GEN_296; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_300 = _GEN_3307 == 10'h241 ? 1'h0 : _GEN_3307 == 10'h241 | (_GEN_3307 == 10'h240 | _GEN_297); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_301 = _GEN_3307 == 10'h242 ? 1'h0 : _GEN_300; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_304 = _GEN_3307 == 10'h243 ? 1'h0 : _GEN_3307 == 10'h243 | (_GEN_3307 == 10'h242 | _GEN_301); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_305 = _GEN_3307 == 10'h244 ? 1'h0 : _GEN_304; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_308 = _GEN_3307 == 10'h245 ? 1'h0 : _GEN_3307 == 10'h245 | (_GEN_3307 == 10'h244 | _GEN_305); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_309 = _GEN_3307 == 10'h246 ? 1'h0 : _GEN_308; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_312 = _GEN_3307 == 10'h247 ? 1'h0 : _GEN_3307 == 10'h247 | (_GEN_3307 == 10'h246 | _GEN_309); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_313 = _GEN_3307 == 10'h248 ? 1'h0 : _GEN_312; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_316 = _GEN_3307 == 10'h249 ? 1'h0 : _GEN_3307 == 10'h249 | (_GEN_3307 == 10'h248 | _GEN_313); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_317 = i == 8'h0 ? 1'h0 : buffer_6; // @[lut_mem_online.scala 210:19 235:34 239:30]
  wire  _GEN_318 = i == 8'h1 ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_319 = i == 8'h8 ? 1'h0 : _GEN_318; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_320 = i == 8'hf ? 1'h0 : _GEN_319; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_321 = i == 8'h11 ? 1'h0 : _GEN_320; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_322 = i == 8'h20 ? 1'h0 : _GEN_321; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_323 = i == 8'h48 ? 1'h0 : _GEN_322; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_324 = _GEN_3306 == 9'h10b ? 1'h0 : _GEN_323; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_325 = _GEN_3306 == 9'h124 ? 1'h0 : _GEN_324; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_326 = _GEN_3307 == 10'h218 ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_328 = _GEN_3307 == 10'h219 ? 1'h0 : _GEN_3307 == 10'h218 | _GEN_326; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_330 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_3307 == 10'h219 | _GEN_328; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_332 = _GEN_3307 == 10'h21b ? 1'h0 : _GEN_3307 == 10'h21a | _GEN_330; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_334 = _GEN_3307 == 10'h21c ? 1'h0 : _GEN_3307 == 10'h21b | _GEN_332; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_336 = _GEN_3307 == 10'h21d ? 1'h0 : _GEN_3307 == 10'h21c | _GEN_334; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_338 = _GEN_3307 == 10'h21e ? 1'h0 : _GEN_3307 == 10'h21d | _GEN_336; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_340 = _GEN_3307 == 10'h21f ? 1'h0 : _GEN_3307 == 10'h21e | _GEN_338; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_342 = _GEN_3307 == 10'h220 ? 1'h0 : _GEN_3307 == 10'h21f | _GEN_340; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_344 = _GEN_3307 == 10'h221 ? 1'h0 : _GEN_3307 == 10'h220 | _GEN_342; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_346 = _GEN_3307 == 10'h222 ? 1'h0 : _GEN_3307 == 10'h221 | _GEN_344; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_348 = _GEN_3307 == 10'h223 ? 1'h0 : _GEN_3307 == 10'h222 | _GEN_346; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_350 = _GEN_3307 == 10'h224 ? 1'h0 : _GEN_3307 == 10'h223 | _GEN_348; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_352 = _GEN_3307 == 10'h225 ? 1'h0 : _GEN_3307 == 10'h224 | _GEN_350; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_354 = _GEN_3307 == 10'h226 ? 1'h0 : _GEN_3307 == 10'h225 | _GEN_352; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_356 = _GEN_3307 == 10'h227 ? 1'h0 : _GEN_3307 == 10'h226 | _GEN_354; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_358 = _GEN_3307 == 10'h228 ? 1'h0 : _GEN_3307 == 10'h227 | _GEN_356; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_360 = _GEN_3307 == 10'h229 ? 1'h0 : _GEN_3307 == 10'h228 | _GEN_358; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_362 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_3307 == 10'h229 | _GEN_360; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_364 = _GEN_3307 == 10'h22b ? 1'h0 : _GEN_3307 == 10'h22a | _GEN_362; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_366 = _GEN_3307 == 10'h22c ? 1'h0 : _GEN_3307 == 10'h22b | _GEN_364; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_368 = _GEN_3307 == 10'h22d ? 1'h0 : _GEN_3307 == 10'h22c | _GEN_366; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_370 = _GEN_3307 == 10'h22e ? 1'h0 : _GEN_3307 == 10'h22d | _GEN_368; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_372 = _GEN_3307 == 10'h22f ? 1'h0 : _GEN_3307 == 10'h22e | _GEN_370; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_374 = _GEN_3307 == 10'h230 ? 1'h0 : _GEN_3307 == 10'h22f | _GEN_372; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_376 = _GEN_3307 == 10'h231 ? 1'h0 : _GEN_3307 == 10'h230 | _GEN_374; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_378 = _GEN_3307 == 10'h232 ? 1'h0 : _GEN_3307 == 10'h231 | _GEN_376; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_380 = _GEN_3307 == 10'h233 ? 1'h0 : _GEN_3307 == 10'h232 | _GEN_378; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_382 = _GEN_3307 == 10'h234 ? 1'h0 : _GEN_3307 == 10'h233 | _GEN_380; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_384 = _GEN_3307 == 10'h235 ? 1'h0 : _GEN_3307 == 10'h234 | _GEN_382; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_386 = _GEN_3307 == 10'h236 ? 1'h0 : _GEN_3307 == 10'h235 | _GEN_384; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_388 = _GEN_3307 == 10'h237 ? 1'h0 : _GEN_3307 == 10'h236 | _GEN_386; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_390 = _GEN_3307 == 10'h238 ? 1'h0 : _GEN_3307 == 10'h237 | _GEN_388; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_392 = _GEN_3307 == 10'h239 ? 1'h0 : _GEN_3307 == 10'h238 | _GEN_390; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_394 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_3307 == 10'h239 | _GEN_392; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_396 = _GEN_3307 == 10'h23b ? 1'h0 : _GEN_3307 == 10'h23a | _GEN_394; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_398 = _GEN_3307 == 10'h23c ? 1'h0 : _GEN_3307 == 10'h23b | _GEN_396; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_400 = _GEN_3307 == 10'h23d ? 1'h0 : _GEN_3307 == 10'h23c | _GEN_398; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_402 = _GEN_3307 == 10'h23e ? 1'h0 : _GEN_3307 == 10'h23d | _GEN_400; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_404 = _GEN_3307 == 10'h23f ? 1'h0 : _GEN_3307 == 10'h23e | _GEN_402; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_406 = _GEN_3307 == 10'h240 ? 1'h0 : _GEN_3307 == 10'h23f | _GEN_404; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_408 = _GEN_3307 == 10'h241 ? 1'h0 : _GEN_3307 == 10'h240 | _GEN_406; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_410 = _GEN_3307 == 10'h242 ? 1'h0 : _GEN_3307 == 10'h241 | _GEN_408; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_412 = _GEN_3307 == 10'h243 ? 1'h0 : _GEN_3307 == 10'h242 | _GEN_410; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_414 = _GEN_3307 == 10'h244 ? 1'h0 : _GEN_3307 == 10'h243 | _GEN_412; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_416 = _GEN_3307 == 10'h245 ? 1'h0 : _GEN_3307 == 10'h244 | _GEN_414; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_418 = _GEN_3307 == 10'h246 ? 1'h0 : _GEN_3307 == 10'h245 | _GEN_416; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_420 = _GEN_3307 == 10'h247 ? 1'h0 : _GEN_3307 == 10'h246 | _GEN_418; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_422 = _GEN_3307 == 10'h248 ? 1'h0 : _GEN_3307 == 10'h247 | _GEN_420; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_424 = _GEN_3307 == 10'h249 ? 1'h0 : _GEN_3307 == 10'h248 | _GEN_422; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_426 = i == 8'h0 ? 1'h0 : _GEN_10; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_427 = i == 8'h1 ? 1'h0 : _GEN_426; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_428 = i == 8'h7 ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_430 = i == 8'h10 ? 1'h0 : i == 8'h8 | _GEN_428; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_432 = i == 8'h22 ? 1'h0 : i == 8'h12 | _GEN_430; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_433 = i == 8'h26 ? 1'h0 : _GEN_432; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_438 = _GEN_3306 == 9'h11b ? 1'h0 : i == 8'h9c | (i == 8'h8d | (i == 8'h4d | (i == 8'h46 | _GEN_433))); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_440 = _GEN_3306 == 9'h13a ? 1'h0 : _GEN_3306 == 9'h11b | _GEN_438; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_442 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_3307 == 10'h275 | _GEN_440; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_443 = i == 8'h0 ? 1'h0 : _GEN_32; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_444 = i == 8'h4 ? 1'h0 : _GEN_443; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_445 = i == 8'h7 ? 1'h0 : _GEN_444; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_446 = i == 8'h9 ? 1'h0 : _GEN_445; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_448 = i == 8'h13 ? 1'h0 : i == 8'h11 | _GEN_446; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_449 = i == 8'h21 ? 1'h0 : _GEN_448; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_451 = i == 8'h23 ? 1'h0 : i == 8'h22 | _GEN_449; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_452 = i == 8'h25 ? 1'h0 : _GEN_451; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_454 = i == 8'h27 ? 1'h0 : i == 8'h26 | _GEN_452; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_456 = i == 8'h46 ? 1'h0 : i == 8'h44 | _GEN_454; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_459 = i == 8'h4d ? 1'h0 : i == 8'h4b | (i == 8'h48 | _GEN_456); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_462 = i == 8'h8d ? 1'h0 : i == 8'h89 | (i == 8'h4f | _GEN_459); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_465 = i == 8'h9c ? 1'h0 : i == 8'h98 | (i == 8'h91 | _GEN_462); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_467 = _GEN_3306 == 9'h113 ? 1'h0 : i == 8'ha0 | _GEN_465; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_470 = _GEN_3306 == 9'h11b ? 1'h0 : _GEN_3306 == 9'h11b | (_GEN_3306 == 9'h113 | _GEN_467); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_471 = _GEN_3306 == 9'h123 ? 1'h0 : _GEN_470; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_473 = _GEN_3306 == 9'h132 ? 1'h0 : _GEN_3306 == 9'h123 | _GEN_471; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_475 = _GEN_3306 == 9'h142 ? 1'h0 : _GEN_3306 == 9'h13a | _GEN_473; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_477 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_3307 == 10'h265 | _GEN_475; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_478 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_477; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_481 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_3307 == 10'h285 | (_GEN_3307 == 10'h275 | _GEN_478); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_482 = i == 8'h0 ? 1'h0 : _GEN_69; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_483 = i == 8'h4 ? 1'h0 : _GEN_482; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_484 = i == 8'h7 ? 1'h0 : _GEN_483; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_485 = i == 8'h9 ? 1'h0 : _GEN_484; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_486 = i == 8'h11 ? 1'h0 : _GEN_485; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_487 = i == 8'h13 ? 1'h0 : _GEN_486; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_489 = i == 8'h44 ? 1'h0 : i == 8'h43 | _GEN_487; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_491 = i == 8'h46 ? 1'h0 : i == 8'h45 | _GEN_489; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_493 = i == 8'h48 ? 1'h0 : i == 8'h47 | _GEN_491; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_494 = i == 8'h4b ? 1'h0 : _GEN_493; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_496 = i == 8'h4d ? 1'h0 : i == 8'h4c | _GEN_494; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_498 = i == 8'h4f ? 1'h0 : i == 8'h4e | _GEN_496; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_501 = i == 8'h89 ? 1'h0 : i == 8'h87 | (i == 8'h50 | _GEN_498); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_503 = i == 8'h8d ? 1'h0 : i == 8'h8b | _GEN_501; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_505 = i == 8'h91 ? 1'h0 : i == 8'h8f | _GEN_503; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_506 = i == 8'h98 ? 1'h0 : _GEN_505; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_508 = i == 8'h9c ? 1'h0 : i == 8'h9a | _GEN_506; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_510 = i == 8'ha0 ? 1'h0 : i == 8'h9e | _GEN_508; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_512 = _GEN_3306 == 9'h10f ? 1'h0 : i == 8'ha2 | _GEN_510; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_515 = _GEN_3306 == 9'h113 ? 1'h0 : _GEN_3306 == 9'h113 | (_GEN_3306 == 9'h10f | _GEN_512); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_516 = _GEN_3306 == 9'h117 ? 1'h0 : _GEN_515; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_519 = _GEN_3306 == 9'h11b ? 1'h0 : _GEN_3306 == 9'h11b | (_GEN_3306 == 9'h117 | _GEN_516); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_520 = _GEN_3306 == 9'h11f ? 1'h0 : _GEN_519; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_523 = _GEN_3306 == 9'h123 ? 1'h0 : _GEN_3306 == 9'h123 | (_GEN_3306 == 9'h11f | _GEN_520); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_525 = _GEN_3306 == 9'h136 ? 1'h0 : _GEN_3306 == 9'h132 | _GEN_523; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_527 = _GEN_3306 == 9'h13e ? 1'h0 : _GEN_3306 == 9'h13a | _GEN_525; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_529 = _GEN_3306 == 9'h146 ? 1'h0 : _GEN_3306 == 9'h142 | _GEN_527; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_530 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_529; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_533 = _GEN_3307 == 10'h26d ? 1'h0 : _GEN_3307 == 10'h26d | (_GEN_3307 == 10'h265 | _GEN_530); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_534 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_533; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_537 = _GEN_3307 == 10'h27d ? 1'h0 : _GEN_3307 == 10'h27d | (_GEN_3307 == 10'h275 | _GEN_534); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_538 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_541 = _GEN_3307 == 10'h28d ? 1'h0 : _GEN_3307 == 10'h28d | (_GEN_3307 == 10'h285 | _GEN_538); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_542 = i == 8'h0 ? 1'h0 : _GEN_124; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_543 = i == 8'h4 ? 1'h0 : _GEN_542; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_544 = i == 8'h9 ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_545 = i == 8'hf ? 1'h0 : _GEN_544; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_546 = i == 8'h11 ? 1'h0 : _GEN_545; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_547 = i == 8'h20 ? 1'h0 : _GEN_546; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_548 = i == 8'h28 ? 1'h0 : _GEN_547; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_549 = i == 8'h42 ? 1'h0 : _GEN_548; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_550 = i == 8'h48 ? 1'h0 : _GEN_549; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_551 = i == 8'h4b ? 1'h0 : _GEN_550; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_552 = i == 8'h51 ? 1'h0 : _GEN_551; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_554 = i == 8'h87 ? 1'h0 : i == 8'h86 | _GEN_552; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_556 = i == 8'h89 ? 1'h0 : i == 8'h88 | _GEN_554; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_558 = i == 8'h8b ? 1'h0 : i == 8'h8a | _GEN_556; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_560 = i == 8'h8d ? 1'h0 : i == 8'h8c | _GEN_558; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_562 = i == 8'h8f ? 1'h0 : i == 8'h8e | _GEN_560; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_564 = i == 8'h91 ? 1'h0 : i == 8'h90 | _GEN_562; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_565 = i == 8'h98 ? 1'h0 : _GEN_564; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_567 = i == 8'h9a ? 1'h0 : i == 8'h99 | _GEN_565; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_569 = i == 8'h9c ? 1'h0 : i == 8'h9b | _GEN_567; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_571 = i == 8'h9e ? 1'h0 : i == 8'h9d | _GEN_569; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_573 = i == 8'ha0 ? 1'h0 : i == 8'h9f | _GEN_571; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_575 = i == 8'ha2 ? 1'h0 : i == 8'ha1 | _GEN_573; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_577 = _GEN_3306 == 9'h10d ? 1'h0 : i == 8'ha3 | _GEN_575; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_580 = _GEN_3306 == 9'h10f ? 1'h0 : _GEN_3306 == 9'h10f | (_GEN_3306 == 9'h10d | _GEN_577); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_581 = _GEN_3306 == 9'h111 ? 1'h0 : _GEN_580; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_584 = _GEN_3306 == 9'h113 ? 1'h0 : _GEN_3306 == 9'h113 | (_GEN_3306 == 9'h111 | _GEN_581); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_585 = _GEN_3306 == 9'h115 ? 1'h0 : _GEN_584; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_588 = _GEN_3306 == 9'h117 ? 1'h0 : _GEN_3306 == 9'h117 | (_GEN_3306 == 9'h115 | _GEN_585); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_589 = _GEN_3306 == 9'h119 ? 1'h0 : _GEN_588; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_592 = _GEN_3306 == 9'h11b ? 1'h0 : _GEN_3306 == 9'h11b | (_GEN_3306 == 9'h119 | _GEN_589); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_593 = _GEN_3306 == 9'h11d ? 1'h0 : _GEN_592; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_596 = _GEN_3306 == 9'h11f ? 1'h0 : _GEN_3306 == 9'h11f | (_GEN_3306 == 9'h11d | _GEN_593); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_597 = _GEN_3306 == 9'h121 ? 1'h0 : _GEN_596; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_600 = _GEN_3306 == 9'h123 ? 1'h0 : _GEN_3306 == 9'h123 | (_GEN_3306 == 9'h121 | _GEN_597); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_602 = _GEN_3306 == 9'h134 ? 1'h0 : _GEN_3306 == 9'h132 | _GEN_600; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_604 = _GEN_3306 == 9'h138 ? 1'h0 : _GEN_3306 == 9'h136 | _GEN_602; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_606 = _GEN_3306 == 9'h13c ? 1'h0 : _GEN_3306 == 9'h13a | _GEN_604; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_608 = _GEN_3306 == 9'h140 ? 1'h0 : _GEN_3306 == 9'h13e | _GEN_606; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_610 = _GEN_3306 == 9'h144 ? 1'h0 : _GEN_3306 == 9'h142 | _GEN_608; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_612 = _GEN_3306 == 9'h148 ? 1'h0 : _GEN_3306 == 9'h146 | _GEN_610; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_613 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_612; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_616 = _GEN_3307 == 10'h269 ? 1'h0 : _GEN_3307 == 10'h269 | (_GEN_3307 == 10'h265 | _GEN_613); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_617 = _GEN_3307 == 10'h26d ? 1'h0 : _GEN_616; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_620 = _GEN_3307 == 10'h271 ? 1'h0 : _GEN_3307 == 10'h271 | (_GEN_3307 == 10'h26d | _GEN_617); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_621 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_620; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_624 = _GEN_3307 == 10'h279 ? 1'h0 : _GEN_3307 == 10'h279 | (_GEN_3307 == 10'h275 | _GEN_621); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_625 = _GEN_3307 == 10'h27d ? 1'h0 : _GEN_624; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_628 = _GEN_3307 == 10'h281 ? 1'h0 : _GEN_3307 == 10'h281 | (_GEN_3307 == 10'h27d | _GEN_625); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_629 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_628; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_632 = _GEN_3307 == 10'h289 ? 1'h0 : _GEN_3307 == 10'h289 | (_GEN_3307 == 10'h285 | _GEN_629); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_633 = _GEN_3307 == 10'h28d ? 1'h0 : _GEN_632; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_636 = _GEN_3307 == 10'h291 ? 1'h0 : _GEN_3307 == 10'h291 | (_GEN_3307 == 10'h28d | _GEN_633); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_637 = i == 8'h0 ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_638 = i == 8'h4 ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_639 = i == 8'h9 ? 1'h0 : _GEN_638; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_640 = i == 8'hf ? 1'h0 : _GEN_639; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_642 = i == 8'h20 ? 1'h0 : i == 8'h11 | _GEN_640; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_643 = i == 8'h28 ? 1'h0 : _GEN_642; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_646 = i == 8'h85 ? 1'h0 : i == 8'h4b | (i == 8'h48 | _GEN_643); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_647 = i == 8'ha4 ? 1'h0 : _GEN_646; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_648 = _GEN_3306 == 9'h10c ? 1'h0 : _GEN_647; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_651 = _GEN_3306 == 9'h10d ? 1'h0 : _GEN_3306 == 9'h10d | (_GEN_3306 == 9'h10c | _GEN_648); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_652 = _GEN_3306 == 9'h10e ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_655 = _GEN_3306 == 9'h10f ? 1'h0 : _GEN_3306 == 9'h10f | (_GEN_3306 == 9'h10e | _GEN_652); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_656 = _GEN_3306 == 9'h110 ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_659 = _GEN_3306 == 9'h111 ? 1'h0 : _GEN_3306 == 9'h111 | (_GEN_3306 == 9'h110 | _GEN_656); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_660 = _GEN_3306 == 9'h112 ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_663 = _GEN_3306 == 9'h113 ? 1'h0 : _GEN_3306 == 9'h113 | (_GEN_3306 == 9'h112 | _GEN_660); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_664 = _GEN_3306 == 9'h114 ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_667 = _GEN_3306 == 9'h115 ? 1'h0 : _GEN_3306 == 9'h115 | (_GEN_3306 == 9'h114 | _GEN_664); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_668 = _GEN_3306 == 9'h116 ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_671 = _GEN_3306 == 9'h117 ? 1'h0 : _GEN_3306 == 9'h117 | (_GEN_3306 == 9'h116 | _GEN_668); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_672 = _GEN_3306 == 9'h118 ? 1'h0 : _GEN_671; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_675 = _GEN_3306 == 9'h119 ? 1'h0 : _GEN_3306 == 9'h119 | (_GEN_3306 == 9'h118 | _GEN_672); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_676 = _GEN_3306 == 9'h11a ? 1'h0 : _GEN_675; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_679 = _GEN_3306 == 9'h11b ? 1'h0 : _GEN_3306 == 9'h11b | (_GEN_3306 == 9'h11a | _GEN_676); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_680 = _GEN_3306 == 9'h11c ? 1'h0 : _GEN_679; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_683 = _GEN_3306 == 9'h11d ? 1'h0 : _GEN_3306 == 9'h11d | (_GEN_3306 == 9'h11c | _GEN_680); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_684 = _GEN_3306 == 9'h11e ? 1'h0 : _GEN_683; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_687 = _GEN_3306 == 9'h11f ? 1'h0 : _GEN_3306 == 9'h11f | (_GEN_3306 == 9'h11e | _GEN_684); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_688 = _GEN_3306 == 9'h120 ? 1'h0 : _GEN_687; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_691 = _GEN_3306 == 9'h121 ? 1'h0 : _GEN_3306 == 9'h121 | (_GEN_3306 == 9'h120 | _GEN_688); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_692 = _GEN_3306 == 9'h122 ? 1'h0 : _GEN_691; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_695 = _GEN_3306 == 9'h123 ? 1'h0 : _GEN_3306 == 9'h123 | (_GEN_3306 == 9'h122 | _GEN_692); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_696 = _GEN_3306 == 9'h124 ? 1'h0 : _GEN_695; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_698 = _GEN_3306 == 9'h131 ? 1'h0 : _GEN_3306 == 9'h124 | _GEN_696; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_700 = _GEN_3306 == 9'h133 ? 1'h0 : _GEN_3306 == 9'h132 | _GEN_698; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_702 = _GEN_3306 == 9'h135 ? 1'h0 : _GEN_3306 == 9'h134 | _GEN_700; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_704 = _GEN_3306 == 9'h137 ? 1'h0 : _GEN_3306 == 9'h136 | _GEN_702; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_706 = _GEN_3306 == 9'h139 ? 1'h0 : _GEN_3306 == 9'h138 | _GEN_704; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_708 = _GEN_3306 == 9'h13b ? 1'h0 : _GEN_3306 == 9'h13a | _GEN_706; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_710 = _GEN_3306 == 9'h13d ? 1'h0 : _GEN_3306 == 9'h13c | _GEN_708; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_712 = _GEN_3306 == 9'h13f ? 1'h0 : _GEN_3306 == 9'h13e | _GEN_710; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_714 = _GEN_3306 == 9'h141 ? 1'h0 : _GEN_3306 == 9'h140 | _GEN_712; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_716 = _GEN_3306 == 9'h143 ? 1'h0 : _GEN_3306 == 9'h142 | _GEN_714; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_718 = _GEN_3306 == 9'h145 ? 1'h0 : _GEN_3306 == 9'h144 | _GEN_716; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_720 = _GEN_3306 == 9'h147 ? 1'h0 : _GEN_3306 == 9'h146 | _GEN_718; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_722 = _GEN_3306 == 9'h149 ? 1'h0 : _GEN_3306 == 9'h148 | _GEN_720; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_724 = _GEN_3307 == 10'h263 ? 1'h0 : _GEN_3307 == 10'h263 | _GEN_722; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_725 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_724; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_728 = _GEN_3307 == 10'h267 ? 1'h0 : _GEN_3307 == 10'h267 | (_GEN_3307 == 10'h265 | _GEN_725); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_729 = _GEN_3307 == 10'h269 ? 1'h0 : _GEN_728; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_732 = _GEN_3307 == 10'h26b ? 1'h0 : _GEN_3307 == 10'h26b | (_GEN_3307 == 10'h269 | _GEN_729); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_733 = _GEN_3307 == 10'h26d ? 1'h0 : _GEN_732; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_736 = _GEN_3307 == 10'h26f ? 1'h0 : _GEN_3307 == 10'h26f | (_GEN_3307 == 10'h26d | _GEN_733); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_737 = _GEN_3307 == 10'h271 ? 1'h0 : _GEN_736; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_740 = _GEN_3307 == 10'h273 ? 1'h0 : _GEN_3307 == 10'h273 | (_GEN_3307 == 10'h271 | _GEN_737); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_741 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_740; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_744 = _GEN_3307 == 10'h277 ? 1'h0 : _GEN_3307 == 10'h277 | (_GEN_3307 == 10'h275 | _GEN_741); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_745 = _GEN_3307 == 10'h279 ? 1'h0 : _GEN_744; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_748 = _GEN_3307 == 10'h27b ? 1'h0 : _GEN_3307 == 10'h27b | (_GEN_3307 == 10'h279 | _GEN_745); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_749 = _GEN_3307 == 10'h27d ? 1'h0 : _GEN_748; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_752 = _GEN_3307 == 10'h27f ? 1'h0 : _GEN_3307 == 10'h27f | (_GEN_3307 == 10'h27d | _GEN_749); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_753 = _GEN_3307 == 10'h281 ? 1'h0 : _GEN_752; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_756 = _GEN_3307 == 10'h283 ? 1'h0 : _GEN_3307 == 10'h283 | (_GEN_3307 == 10'h281 | _GEN_753); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_757 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_756; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_760 = _GEN_3307 == 10'h287 ? 1'h0 : _GEN_3307 == 10'h287 | (_GEN_3307 == 10'h285 | _GEN_757); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_761 = _GEN_3307 == 10'h289 ? 1'h0 : _GEN_760; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_764 = _GEN_3307 == 10'h28b ? 1'h0 : _GEN_3307 == 10'h28b | (_GEN_3307 == 10'h289 | _GEN_761); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_765 = _GEN_3307 == 10'h28d ? 1'h0 : _GEN_764; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_768 = _GEN_3307 == 10'h28f ? 1'h0 : _GEN_3307 == 10'h28f | (_GEN_3307 == 10'h28d | _GEN_765); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_769 = _GEN_3307 == 10'h291 ? 1'h0 : _GEN_768; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_772 = _GEN_3307 == 10'h293 ? 1'h0 : _GEN_3307 == 10'h293 | (_GEN_3307 == 10'h291 | _GEN_769); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_773 = i == 8'h0 ? 1'h0 : _GEN_316; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_774 = i == 8'h4 ? 1'h0 : _GEN_773; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_775 = i == 8'h9 ? 1'h0 : _GEN_774; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_776 = i == 8'hf ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_777 = i == 8'h11 ? 1'h0 : _GEN_776; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_778 = i == 8'h20 ? 1'h0 : _GEN_777; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_779 = i == 8'h28 ? 1'h0 : _GEN_778; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_780 = i == 8'h48 ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_781 = i == 8'h4b ? 1'h0 : _GEN_780; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_782 = i == 8'h85 ? 1'h0 : _GEN_781; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_783 = i == 8'ha4 ? 1'h0 : _GEN_782; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_785 = _GEN_3306 == 9'h10c ? 1'h0 : _GEN_3306 == 9'h10c | _GEN_783; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_787 = _GEN_3306 == 9'h10d ? 1'h0 : _GEN_3306 == 9'h10d | _GEN_785; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_789 = _GEN_3306 == 9'h10e ? 1'h0 : _GEN_3306 == 9'h10e | _GEN_787; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_791 = _GEN_3306 == 9'h10f ? 1'h0 : _GEN_3306 == 9'h10f | _GEN_789; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_793 = _GEN_3306 == 9'h110 ? 1'h0 : _GEN_3306 == 9'h110 | _GEN_791; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_795 = _GEN_3306 == 9'h111 ? 1'h0 : _GEN_3306 == 9'h111 | _GEN_793; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_797 = _GEN_3306 == 9'h112 ? 1'h0 : _GEN_3306 == 9'h112 | _GEN_795; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_799 = _GEN_3306 == 9'h113 ? 1'h0 : _GEN_3306 == 9'h113 | _GEN_797; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_801 = _GEN_3306 == 9'h114 ? 1'h0 : _GEN_3306 == 9'h114 | _GEN_799; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_803 = _GEN_3306 == 9'h115 ? 1'h0 : _GEN_3306 == 9'h115 | _GEN_801; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_805 = _GEN_3306 == 9'h116 ? 1'h0 : _GEN_3306 == 9'h116 | _GEN_803; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_807 = _GEN_3306 == 9'h117 ? 1'h0 : _GEN_3306 == 9'h117 | _GEN_805; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_809 = _GEN_3306 == 9'h118 ? 1'h0 : _GEN_3306 == 9'h118 | _GEN_807; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_811 = _GEN_3306 == 9'h119 ? 1'h0 : _GEN_3306 == 9'h119 | _GEN_809; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_813 = _GEN_3306 == 9'h11a ? 1'h0 : _GEN_3306 == 9'h11a | _GEN_811; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_815 = _GEN_3306 == 9'h11b ? 1'h0 : _GEN_3306 == 9'h11b | _GEN_813; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_817 = _GEN_3306 == 9'h11c ? 1'h0 : _GEN_3306 == 9'h11c | _GEN_815; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_819 = _GEN_3306 == 9'h11d ? 1'h0 : _GEN_3306 == 9'h11d | _GEN_817; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_821 = _GEN_3306 == 9'h11e ? 1'h0 : _GEN_3306 == 9'h11e | _GEN_819; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_823 = _GEN_3306 == 9'h11f ? 1'h0 : _GEN_3306 == 9'h11f | _GEN_821; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_825 = _GEN_3306 == 9'h120 ? 1'h0 : _GEN_3306 == 9'h120 | _GEN_823; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_827 = _GEN_3306 == 9'h121 ? 1'h0 : _GEN_3306 == 9'h121 | _GEN_825; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_829 = _GEN_3306 == 9'h122 ? 1'h0 : _GEN_3306 == 9'h122 | _GEN_827; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_831 = _GEN_3306 == 9'h123 ? 1'h0 : _GEN_3306 == 9'h123 | _GEN_829; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_833 = _GEN_3306 == 9'h124 ? 1'h0 : _GEN_3306 == 9'h124 | _GEN_831; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_834 = _GEN_3307 == 10'h263 ? 1'h0 : _GEN_833; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_837 = _GEN_3307 == 10'h264 ? 1'h0 : _GEN_3307 == 10'h264 | (_GEN_3307 == 10'h263 | _GEN_834); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_838 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_837; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_841 = _GEN_3307 == 10'h266 ? 1'h0 : _GEN_3307 == 10'h266 | (_GEN_3307 == 10'h265 | _GEN_838); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_842 = _GEN_3307 == 10'h267 ? 1'h0 : _GEN_841; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_845 = _GEN_3307 == 10'h268 ? 1'h0 : _GEN_3307 == 10'h268 | (_GEN_3307 == 10'h267 | _GEN_842); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_846 = _GEN_3307 == 10'h269 ? 1'h0 : _GEN_845; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_849 = _GEN_3307 == 10'h26a ? 1'h0 : _GEN_3307 == 10'h26a | (_GEN_3307 == 10'h269 | _GEN_846); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_850 = _GEN_3307 == 10'h26b ? 1'h0 : _GEN_849; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_853 = _GEN_3307 == 10'h26c ? 1'h0 : _GEN_3307 == 10'h26c | (_GEN_3307 == 10'h26b | _GEN_850); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_854 = _GEN_3307 == 10'h26d ? 1'h0 : _GEN_853; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_857 = _GEN_3307 == 10'h26e ? 1'h0 : _GEN_3307 == 10'h26e | (_GEN_3307 == 10'h26d | _GEN_854); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_858 = _GEN_3307 == 10'h26f ? 1'h0 : _GEN_857; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_861 = _GEN_3307 == 10'h270 ? 1'h0 : _GEN_3307 == 10'h270 | (_GEN_3307 == 10'h26f | _GEN_858); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_862 = _GEN_3307 == 10'h271 ? 1'h0 : _GEN_861; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_865 = _GEN_3307 == 10'h272 ? 1'h0 : _GEN_3307 == 10'h272 | (_GEN_3307 == 10'h271 | _GEN_862); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_866 = _GEN_3307 == 10'h273 ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_869 = _GEN_3307 == 10'h274 ? 1'h0 : _GEN_3307 == 10'h274 | (_GEN_3307 == 10'h273 | _GEN_866); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_870 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_869; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_873 = _GEN_3307 == 10'h276 ? 1'h0 : _GEN_3307 == 10'h276 | (_GEN_3307 == 10'h275 | _GEN_870); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_874 = _GEN_3307 == 10'h277 ? 1'h0 : _GEN_873; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_877 = _GEN_3307 == 10'h278 ? 1'h0 : _GEN_3307 == 10'h278 | (_GEN_3307 == 10'h277 | _GEN_874); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_878 = _GEN_3307 == 10'h279 ? 1'h0 : _GEN_877; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_881 = _GEN_3307 == 10'h27a ? 1'h0 : _GEN_3307 == 10'h27a | (_GEN_3307 == 10'h279 | _GEN_878); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_882 = _GEN_3307 == 10'h27b ? 1'h0 : _GEN_881; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_885 = _GEN_3307 == 10'h27c ? 1'h0 : _GEN_3307 == 10'h27c | (_GEN_3307 == 10'h27b | _GEN_882); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_886 = _GEN_3307 == 10'h27d ? 1'h0 : _GEN_885; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_889 = _GEN_3307 == 10'h27e ? 1'h0 : _GEN_3307 == 10'h27e | (_GEN_3307 == 10'h27d | _GEN_886); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_890 = _GEN_3307 == 10'h27f ? 1'h0 : _GEN_889; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_893 = _GEN_3307 == 10'h280 ? 1'h0 : _GEN_3307 == 10'h280 | (_GEN_3307 == 10'h27f | _GEN_890); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_894 = _GEN_3307 == 10'h281 ? 1'h0 : _GEN_893; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_897 = _GEN_3307 == 10'h282 ? 1'h0 : _GEN_3307 == 10'h282 | (_GEN_3307 == 10'h281 | _GEN_894); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_898 = _GEN_3307 == 10'h283 ? 1'h0 : _GEN_897; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_901 = _GEN_3307 == 10'h284 ? 1'h0 : _GEN_3307 == 10'h284 | (_GEN_3307 == 10'h283 | _GEN_898); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_902 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_901; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_905 = _GEN_3307 == 10'h286 ? 1'h0 : _GEN_3307 == 10'h286 | (_GEN_3307 == 10'h285 | _GEN_902); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_906 = _GEN_3307 == 10'h287 ? 1'h0 : _GEN_905; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_909 = _GEN_3307 == 10'h288 ? 1'h0 : _GEN_3307 == 10'h288 | (_GEN_3307 == 10'h287 | _GEN_906); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_910 = _GEN_3307 == 10'h289 ? 1'h0 : _GEN_909; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_913 = _GEN_3307 == 10'h28a ? 1'h0 : _GEN_3307 == 10'h28a | (_GEN_3307 == 10'h289 | _GEN_910); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_914 = _GEN_3307 == 10'h28b ? 1'h0 : _GEN_913; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_917 = _GEN_3307 == 10'h28c ? 1'h0 : _GEN_3307 == 10'h28c | (_GEN_3307 == 10'h28b | _GEN_914); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_918 = _GEN_3307 == 10'h28d ? 1'h0 : _GEN_917; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_921 = _GEN_3307 == 10'h28e ? 1'h0 : _GEN_3307 == 10'h28e | (_GEN_3307 == 10'h28d | _GEN_918); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_922 = _GEN_3307 == 10'h28f ? 1'h0 : _GEN_921; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_925 = _GEN_3307 == 10'h290 ? 1'h0 : _GEN_3307 == 10'h290 | (_GEN_3307 == 10'h28f | _GEN_922); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_926 = _GEN_3307 == 10'h291 ? 1'h0 : _GEN_925; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_929 = _GEN_3307 == 10'h292 ? 1'h0 : _GEN_3307 == 10'h292 | (_GEN_3307 == 10'h291 | _GEN_926); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_930 = _GEN_3307 == 10'h293 ? 1'h0 : _GEN_929; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_933 = _GEN_3307 == 10'h294 ? 1'h0 : _GEN_3307 == 10'h294 | (_GEN_3307 == 10'h293 | _GEN_930); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_934 = i == 8'h0 ? 1'h0 : _GEN_3307 == 10'h249 | _GEN_424; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_935 = i == 8'h4 ? 1'h0 : _GEN_934; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_936 = i == 8'h9 ? 1'h0 : _GEN_935; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_937 = i == 8'hf ? 1'h0 : _GEN_936; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_938 = i == 8'h11 ? 1'h0 : _GEN_937; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_939 = i == 8'h20 ? 1'h0 : _GEN_938; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_940 = i == 8'h28 ? 1'h0 : _GEN_939; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_941 = i == 8'h48 ? 1'h0 : _GEN_940; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_942 = i == 8'h4b ? 1'h0 : _GEN_941; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_943 = i == 8'ha4 ? 1'h0 : _GEN_942; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_944 = _GEN_3306 == 9'h10b ? 1'h0 : _GEN_943; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_945 = _GEN_3306 == 9'h124 ? 1'h0 : _GEN_944; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_946 = _GEN_3307 == 10'h218 ? 1'h0 : _GEN_945; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_948 = _GEN_3307 == 10'h219 ? 1'h0 : _GEN_3307 == 10'h218 | _GEN_946; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_950 = _GEN_3307 == 10'h21a ? 1'h0 : _GEN_3307 == 10'h219 | _GEN_948; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_952 = _GEN_3307 == 10'h21b ? 1'h0 : _GEN_3307 == 10'h21a | _GEN_950; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_954 = _GEN_3307 == 10'h21c ? 1'h0 : _GEN_3307 == 10'h21b | _GEN_952; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_956 = _GEN_3307 == 10'h21d ? 1'h0 : _GEN_3307 == 10'h21c | _GEN_954; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_958 = _GEN_3307 == 10'h21e ? 1'h0 : _GEN_3307 == 10'h21d | _GEN_956; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_960 = _GEN_3307 == 10'h21f ? 1'h0 : _GEN_3307 == 10'h21e | _GEN_958; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_962 = _GEN_3307 == 10'h220 ? 1'h0 : _GEN_3307 == 10'h21f | _GEN_960; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_964 = _GEN_3307 == 10'h221 ? 1'h0 : _GEN_3307 == 10'h220 | _GEN_962; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_966 = _GEN_3307 == 10'h222 ? 1'h0 : _GEN_3307 == 10'h221 | _GEN_964; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_968 = _GEN_3307 == 10'h223 ? 1'h0 : _GEN_3307 == 10'h222 | _GEN_966; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_970 = _GEN_3307 == 10'h224 ? 1'h0 : _GEN_3307 == 10'h223 | _GEN_968; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_972 = _GEN_3307 == 10'h225 ? 1'h0 : _GEN_3307 == 10'h224 | _GEN_970; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_974 = _GEN_3307 == 10'h226 ? 1'h0 : _GEN_3307 == 10'h225 | _GEN_972; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_976 = _GEN_3307 == 10'h227 ? 1'h0 : _GEN_3307 == 10'h226 | _GEN_974; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_978 = _GEN_3307 == 10'h228 ? 1'h0 : _GEN_3307 == 10'h227 | _GEN_976; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_980 = _GEN_3307 == 10'h229 ? 1'h0 : _GEN_3307 == 10'h228 | _GEN_978; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_982 = _GEN_3307 == 10'h22a ? 1'h0 : _GEN_3307 == 10'h229 | _GEN_980; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_984 = _GEN_3307 == 10'h22b ? 1'h0 : _GEN_3307 == 10'h22a | _GEN_982; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_986 = _GEN_3307 == 10'h22c ? 1'h0 : _GEN_3307 == 10'h22b | _GEN_984; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_988 = _GEN_3307 == 10'h22d ? 1'h0 : _GEN_3307 == 10'h22c | _GEN_986; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_990 = _GEN_3307 == 10'h22e ? 1'h0 : _GEN_3307 == 10'h22d | _GEN_988; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_992 = _GEN_3307 == 10'h22f ? 1'h0 : _GEN_3307 == 10'h22e | _GEN_990; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_994 = _GEN_3307 == 10'h230 ? 1'h0 : _GEN_3307 == 10'h22f | _GEN_992; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_996 = _GEN_3307 == 10'h231 ? 1'h0 : _GEN_3307 == 10'h230 | _GEN_994; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_998 = _GEN_3307 == 10'h232 ? 1'h0 : _GEN_3307 == 10'h231 | _GEN_996; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1000 = _GEN_3307 == 10'h233 ? 1'h0 : _GEN_3307 == 10'h232 | _GEN_998; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1002 = _GEN_3307 == 10'h234 ? 1'h0 : _GEN_3307 == 10'h233 | _GEN_1000; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1004 = _GEN_3307 == 10'h235 ? 1'h0 : _GEN_3307 == 10'h234 | _GEN_1002; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1006 = _GEN_3307 == 10'h236 ? 1'h0 : _GEN_3307 == 10'h235 | _GEN_1004; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1008 = _GEN_3307 == 10'h237 ? 1'h0 : _GEN_3307 == 10'h236 | _GEN_1006; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1010 = _GEN_3307 == 10'h238 ? 1'h0 : _GEN_3307 == 10'h237 | _GEN_1008; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1012 = _GEN_3307 == 10'h239 ? 1'h0 : _GEN_3307 == 10'h238 | _GEN_1010; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1014 = _GEN_3307 == 10'h23a ? 1'h0 : _GEN_3307 == 10'h239 | _GEN_1012; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1016 = _GEN_3307 == 10'h23b ? 1'h0 : _GEN_3307 == 10'h23a | _GEN_1014; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1018 = _GEN_3307 == 10'h23c ? 1'h0 : _GEN_3307 == 10'h23b | _GEN_1016; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1020 = _GEN_3307 == 10'h23d ? 1'h0 : _GEN_3307 == 10'h23c | _GEN_1018; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1022 = _GEN_3307 == 10'h23e ? 1'h0 : _GEN_3307 == 10'h23d | _GEN_1020; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1024 = _GEN_3307 == 10'h23f ? 1'h0 : _GEN_3307 == 10'h23e | _GEN_1022; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1026 = _GEN_3307 == 10'h240 ? 1'h0 : _GEN_3307 == 10'h23f | _GEN_1024; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1028 = _GEN_3307 == 10'h241 ? 1'h0 : _GEN_3307 == 10'h240 | _GEN_1026; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1030 = _GEN_3307 == 10'h242 ? 1'h0 : _GEN_3307 == 10'h241 | _GEN_1028; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1032 = _GEN_3307 == 10'h243 ? 1'h0 : _GEN_3307 == 10'h242 | _GEN_1030; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1034 = _GEN_3307 == 10'h244 ? 1'h0 : _GEN_3307 == 10'h243 | _GEN_1032; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1036 = _GEN_3307 == 10'h245 ? 1'h0 : _GEN_3307 == 10'h244 | _GEN_1034; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1038 = _GEN_3307 == 10'h246 ? 1'h0 : _GEN_3307 == 10'h245 | _GEN_1036; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1040 = _GEN_3307 == 10'h247 ? 1'h0 : _GEN_3307 == 10'h246 | _GEN_1038; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1042 = _GEN_3307 == 10'h248 ? 1'h0 : _GEN_3307 == 10'h247 | _GEN_1040; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1044 = _GEN_3307 == 10'h249 ? 1'h0 : _GEN_3307 == 10'h248 | _GEN_1042; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1046 = _GEN_3307 == 10'h263 ? 1'h0 : _GEN_3307 == 10'h249 | _GEN_1044; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1048 = _GEN_3307 == 10'h264 ? 1'h0 : _GEN_3307 == 10'h263 | _GEN_1046; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1050 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_3307 == 10'h264 | _GEN_1048; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1052 = _GEN_3307 == 10'h266 ? 1'h0 : _GEN_3307 == 10'h265 | _GEN_1050; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1054 = _GEN_3307 == 10'h267 ? 1'h0 : _GEN_3307 == 10'h266 | _GEN_1052; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1056 = _GEN_3307 == 10'h268 ? 1'h0 : _GEN_3307 == 10'h267 | _GEN_1054; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1058 = _GEN_3307 == 10'h269 ? 1'h0 : _GEN_3307 == 10'h268 | _GEN_1056; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1060 = _GEN_3307 == 10'h26a ? 1'h0 : _GEN_3307 == 10'h269 | _GEN_1058; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1062 = _GEN_3307 == 10'h26b ? 1'h0 : _GEN_3307 == 10'h26a | _GEN_1060; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1064 = _GEN_3307 == 10'h26c ? 1'h0 : _GEN_3307 == 10'h26b | _GEN_1062; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1066 = _GEN_3307 == 10'h26d ? 1'h0 : _GEN_3307 == 10'h26c | _GEN_1064; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1068 = _GEN_3307 == 10'h26e ? 1'h0 : _GEN_3307 == 10'h26d | _GEN_1066; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1070 = _GEN_3307 == 10'h26f ? 1'h0 : _GEN_3307 == 10'h26e | _GEN_1068; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1072 = _GEN_3307 == 10'h270 ? 1'h0 : _GEN_3307 == 10'h26f | _GEN_1070; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1074 = _GEN_3307 == 10'h271 ? 1'h0 : _GEN_3307 == 10'h270 | _GEN_1072; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1076 = _GEN_3307 == 10'h272 ? 1'h0 : _GEN_3307 == 10'h271 | _GEN_1074; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1078 = _GEN_3307 == 10'h273 ? 1'h0 : _GEN_3307 == 10'h272 | _GEN_1076; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1080 = _GEN_3307 == 10'h274 ? 1'h0 : _GEN_3307 == 10'h273 | _GEN_1078; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1082 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_3307 == 10'h274 | _GEN_1080; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1084 = _GEN_3307 == 10'h276 ? 1'h0 : _GEN_3307 == 10'h275 | _GEN_1082; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1086 = _GEN_3307 == 10'h277 ? 1'h0 : _GEN_3307 == 10'h276 | _GEN_1084; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1088 = _GEN_3307 == 10'h278 ? 1'h0 : _GEN_3307 == 10'h277 | _GEN_1086; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1090 = _GEN_3307 == 10'h279 ? 1'h0 : _GEN_3307 == 10'h278 | _GEN_1088; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1092 = _GEN_3307 == 10'h27a ? 1'h0 : _GEN_3307 == 10'h279 | _GEN_1090; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1094 = _GEN_3307 == 10'h27b ? 1'h0 : _GEN_3307 == 10'h27a | _GEN_1092; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1096 = _GEN_3307 == 10'h27c ? 1'h0 : _GEN_3307 == 10'h27b | _GEN_1094; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1098 = _GEN_3307 == 10'h27d ? 1'h0 : _GEN_3307 == 10'h27c | _GEN_1096; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1100 = _GEN_3307 == 10'h27e ? 1'h0 : _GEN_3307 == 10'h27d | _GEN_1098; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1102 = _GEN_3307 == 10'h27f ? 1'h0 : _GEN_3307 == 10'h27e | _GEN_1100; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1104 = _GEN_3307 == 10'h280 ? 1'h0 : _GEN_3307 == 10'h27f | _GEN_1102; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1106 = _GEN_3307 == 10'h281 ? 1'h0 : _GEN_3307 == 10'h280 | _GEN_1104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1108 = _GEN_3307 == 10'h282 ? 1'h0 : _GEN_3307 == 10'h281 | _GEN_1106; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1110 = _GEN_3307 == 10'h283 ? 1'h0 : _GEN_3307 == 10'h282 | _GEN_1108; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1112 = _GEN_3307 == 10'h284 ? 1'h0 : _GEN_3307 == 10'h283 | _GEN_1110; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1114 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_3307 == 10'h284 | _GEN_1112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1116 = _GEN_3307 == 10'h286 ? 1'h0 : _GEN_3307 == 10'h285 | _GEN_1114; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1118 = _GEN_3307 == 10'h287 ? 1'h0 : _GEN_3307 == 10'h286 | _GEN_1116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1120 = _GEN_3307 == 10'h288 ? 1'h0 : _GEN_3307 == 10'h287 | _GEN_1118; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1122 = _GEN_3307 == 10'h289 ? 1'h0 : _GEN_3307 == 10'h288 | _GEN_1120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1124 = _GEN_3307 == 10'h28a ? 1'h0 : _GEN_3307 == 10'h289 | _GEN_1122; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1126 = _GEN_3307 == 10'h28b ? 1'h0 : _GEN_3307 == 10'h28a | _GEN_1124; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1128 = _GEN_3307 == 10'h28c ? 1'h0 : _GEN_3307 == 10'h28b | _GEN_1126; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1130 = _GEN_3307 == 10'h28d ? 1'h0 : _GEN_3307 == 10'h28c | _GEN_1128; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1132 = _GEN_3307 == 10'h28e ? 1'h0 : _GEN_3307 == 10'h28d | _GEN_1130; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1134 = _GEN_3307 == 10'h28f ? 1'h0 : _GEN_3307 == 10'h28e | _GEN_1132; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1136 = _GEN_3307 == 10'h290 ? 1'h0 : _GEN_3307 == 10'h28f | _GEN_1134; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1138 = _GEN_3307 == 10'h291 ? 1'h0 : _GEN_3307 == 10'h290 | _GEN_1136; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1140 = _GEN_3307 == 10'h292 ? 1'h0 : _GEN_3307 == 10'h291 | _GEN_1138; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1142 = _GEN_3307 == 10'h293 ? 1'h0 : _GEN_3307 == 10'h292 | _GEN_1140; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1144 = _GEN_3307 == 10'h294 ? 1'h0 : _GEN_3307 == 10'h293 | _GEN_1142; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1146 = i == 8'h0 ? 1'h0 : _GEN_442; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1147 = i == 8'h1 ? 1'h0 : _GEN_1146; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1148 = i == 8'h4 ? 1'h0 : _GEN_1147; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1149 = i == 8'h9 ? 1'h0 : _GEN_1148; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1151 = i == 8'h28 ? 1'h0 : i == 8'h27 | _GEN_1149; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1152 = i == 8'h4f ? 1'h0 : _GEN_1151; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1156 = _GEN_3306 == 9'h14a ? 1'h0 : i == 8'ha4 | (i == 8'h51 | (i == 8'h4f | _GEN_1152)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1158 = _GEN_3307 == 10'h295 ? 1'h0 : _GEN_3307 == 10'h295 | _GEN_1156; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1159 = i == 8'h0 ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1160 = i == 8'h3 ? 1'h0 : _GEN_1159; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1161 = i == 8'h4 ? 1'h0 : _GEN_1160; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1162 = i == 8'h8 ? 1'h0 : _GEN_1161; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1163 = i == 8'h9 ? 1'h0 : _GEN_1162; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1164 = i == 8'h12 ? 1'h0 : _GEN_1163; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1166 = i == 8'h27 ? 1'h0 : i == 8'h26 | _GEN_1164; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1167 = i == 8'h28 ? 1'h0 : _GEN_1166; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1168 = i == 8'h4d ? 1'h0 : _GEN_1167; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1171 = i == 8'h4f ? 1'h0 : i == 8'h4f | (i == 8'h4d | _GEN_1168); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1172 = i == 8'h51 ? 1'h0 : _GEN_1171; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1174 = _GEN_3306 == 9'h14a ? 1'h0 : i == 8'ha4 | _GEN_1172; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1176 = _GEN_3307 == 10'h295 ? 1'h0 : _GEN_3307 == 10'h295 | _GEN_1174; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1177 = i == 8'h0 ? 1'h0 : _GEN_541; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1178 = i == 8'h3 ? 1'h0 : _GEN_1177; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1179 = i == 8'h4 ? 1'h0 : _GEN_1178; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1180 = i == 8'h8 ? 1'h0 : _GEN_1179; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1181 = i == 8'h9 ? 1'h0 : _GEN_1180; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1182 = i == 8'h25 ? 1'h0 : _GEN_1181; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1183 = i == 8'h28 ? 1'h0 : _GEN_1182; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1184 = i == 8'h4c ? 1'h0 : _GEN_1183; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1187 = i == 8'h4d ? 1'h0 : i == 8'h4d | (i == 8'h4c | _GEN_1184); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1188 = i == 8'h4e ? 1'h0 : _GEN_1187; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1191 = i == 8'h4f ? 1'h0 : i == 8'h4f | (i == 8'h4e | _GEN_1188); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1192 = i == 8'h50 ? 1'h0 : _GEN_1191; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1195 = i == 8'h51 ? 1'h0 : i == 8'h51 | (i == 8'h50 | _GEN_1192); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1196 = i == 8'h0 ? 1'h0 : _GEN_636; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1197 = i == 8'h3 ? 1'h0 : _GEN_1196; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1198 = i == 8'h4 ? 1'h0 : _GEN_1197; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1199 = i == 8'h8 ? 1'h0 : _GEN_1198; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1200 = i == 8'h9 ? 1'h0 : _GEN_1199; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1201 = i == 8'h25 ? 1'h0 : _GEN_1200; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1202 = i == 8'h28 ? 1'h0 : _GEN_1201; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1204 = i == 8'h4c ? 1'h0 : i == 8'h4c | _GEN_1202; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1206 = i == 8'h4d ? 1'h0 : i == 8'h4d | _GEN_1204; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1208 = i == 8'h4e ? 1'h0 : i == 8'h4e | _GEN_1206; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1210 = i == 8'h4f ? 1'h0 : i == 8'h4f | _GEN_1208; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1212 = i == 8'h50 ? 1'h0 : i == 8'h50 | _GEN_1210; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1214 = i == 8'h51 ? 1'h0 : i == 8'h51 | _GEN_1212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1215 = i == 8'h0 ? 1'h0 : _GEN_772; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1216 = i == 8'h3 ? 1'h0 : _GEN_1215; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1217 = i == 8'h4 ? 1'h0 : _GEN_1216; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1218 = i == 8'h8 ? 1'h0 : _GEN_1217; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1219 = i == 8'h9 ? 1'h0 : _GEN_1218; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1220 = i == 8'h28 ? 1'h0 : _GEN_1219; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1221 = i == 8'h4b ? 1'h0 : _GEN_1220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1222 = i == 8'h98 ? 1'h0 : _GEN_1221; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1224 = i == 8'h99 ? 1'h0 : i == 8'h98 | _GEN_1222; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1226 = i == 8'h9a ? 1'h0 : i == 8'h99 | _GEN_1224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1228 = i == 8'h9b ? 1'h0 : i == 8'h9a | _GEN_1226; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1230 = i == 8'h9c ? 1'h0 : i == 8'h9b | _GEN_1228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1232 = i == 8'h9d ? 1'h0 : i == 8'h9c | _GEN_1230; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1234 = i == 8'h9e ? 1'h0 : i == 8'h9d | _GEN_1232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1236 = i == 8'h9f ? 1'h0 : i == 8'h9e | _GEN_1234; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1238 = i == 8'ha0 ? 1'h0 : i == 8'h9f | _GEN_1236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1240 = i == 8'ha1 ? 1'h0 : i == 8'ha0 | _GEN_1238; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1242 = i == 8'ha2 ? 1'h0 : i == 8'ha1 | _GEN_1240; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1244 = i == 8'ha3 ? 1'h0 : i == 8'ha2 | _GEN_1242; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1246 = i == 8'ha4 ? 1'h0 : i == 8'ha3 | _GEN_1244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1247 = _GEN_3306 == 9'h14a ? 1'h0 : _GEN_1246; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1249 = _GEN_3307 == 10'h295 ? 1'h0 : _GEN_3307 == 10'h295 | _GEN_1247; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1250 = i == 8'h0 ? 1'h0 : _GEN_933; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1251 = i == 8'h3 ? 1'h0 : _GEN_1250; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1252 = i == 8'h4 ? 1'h0 : _GEN_1251; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1253 = i == 8'h8 ? 1'h0 : _GEN_1252; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1254 = i == 8'h9 ? 1'h0 : _GEN_1253; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1255 = i == 8'h28 ? 1'h0 : _GEN_1254; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1256 = i == 8'h4b ? 1'h0 : _GEN_1255; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1257 = i == 8'ha4 ? 1'h0 : _GEN_1256; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1258 = _GEN_3306 == 9'h131 ? 1'h0 : _GEN_1257; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1260 = _GEN_3306 == 9'h132 ? 1'h0 : _GEN_3306 == 9'h131 | _GEN_1258; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1262 = _GEN_3306 == 9'h133 ? 1'h0 : _GEN_3306 == 9'h132 | _GEN_1260; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1264 = _GEN_3306 == 9'h134 ? 1'h0 : _GEN_3306 == 9'h133 | _GEN_1262; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1266 = _GEN_3306 == 9'h135 ? 1'h0 : _GEN_3306 == 9'h134 | _GEN_1264; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1268 = _GEN_3306 == 9'h136 ? 1'h0 : _GEN_3306 == 9'h135 | _GEN_1266; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1270 = _GEN_3306 == 9'h137 ? 1'h0 : _GEN_3306 == 9'h136 | _GEN_1268; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1272 = _GEN_3306 == 9'h138 ? 1'h0 : _GEN_3306 == 9'h137 | _GEN_1270; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1274 = _GEN_3306 == 9'h139 ? 1'h0 : _GEN_3306 == 9'h138 | _GEN_1272; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1276 = _GEN_3306 == 9'h13a ? 1'h0 : _GEN_3306 == 9'h139 | _GEN_1274; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1278 = _GEN_3306 == 9'h13b ? 1'h0 : _GEN_3306 == 9'h13a | _GEN_1276; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1280 = _GEN_3306 == 9'h13c ? 1'h0 : _GEN_3306 == 9'h13b | _GEN_1278; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1282 = _GEN_3306 == 9'h13d ? 1'h0 : _GEN_3306 == 9'h13c | _GEN_1280; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1284 = _GEN_3306 == 9'h13e ? 1'h0 : _GEN_3306 == 9'h13d | _GEN_1282; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1286 = _GEN_3306 == 9'h13f ? 1'h0 : _GEN_3306 == 9'h13e | _GEN_1284; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1288 = _GEN_3306 == 9'h140 ? 1'h0 : _GEN_3306 == 9'h13f | _GEN_1286; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1290 = _GEN_3306 == 9'h141 ? 1'h0 : _GEN_3306 == 9'h140 | _GEN_1288; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1292 = _GEN_3306 == 9'h142 ? 1'h0 : _GEN_3306 == 9'h141 | _GEN_1290; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1294 = _GEN_3306 == 9'h143 ? 1'h0 : _GEN_3306 == 9'h142 | _GEN_1292; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1296 = _GEN_3306 == 9'h144 ? 1'h0 : _GEN_3306 == 9'h143 | _GEN_1294; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1298 = _GEN_3306 == 9'h145 ? 1'h0 : _GEN_3306 == 9'h144 | _GEN_1296; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1300 = _GEN_3306 == 9'h146 ? 1'h0 : _GEN_3306 == 9'h145 | _GEN_1298; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1302 = _GEN_3306 == 9'h147 ? 1'h0 : _GEN_3306 == 9'h146 | _GEN_1300; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1304 = _GEN_3306 == 9'h148 ? 1'h0 : _GEN_3306 == 9'h147 | _GEN_1302; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1306 = _GEN_3306 == 9'h149 ? 1'h0 : _GEN_3306 == 9'h148 | _GEN_1304; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1308 = i == 8'h0 ? 1'h0 : _GEN_3307 == 10'h294 | _GEN_1144; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1309 = i == 8'h3 ? 1'h0 : _GEN_1308; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1310 = i == 8'h4 ? 1'h0 : _GEN_1309; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1311 = i == 8'h8 ? 1'h0 : _GEN_1310; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1312 = i == 8'h9 ? 1'h0 : _GEN_1311; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1313 = i == 8'h28 ? 1'h0 : _GEN_1312; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1314 = i == 8'h4b ? 1'h0 : _GEN_1313; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1315 = i == 8'ha4 ? 1'h0 : _GEN_1314; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1316 = _GEN_3307 == 10'h263 ? 1'h0 : _GEN_1315; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1318 = _GEN_3307 == 10'h264 ? 1'h0 : _GEN_3307 == 10'h263 | _GEN_1316; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1320 = _GEN_3307 == 10'h265 ? 1'h0 : _GEN_3307 == 10'h264 | _GEN_1318; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1322 = _GEN_3307 == 10'h266 ? 1'h0 : _GEN_3307 == 10'h265 | _GEN_1320; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1324 = _GEN_3307 == 10'h267 ? 1'h0 : _GEN_3307 == 10'h266 | _GEN_1322; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1326 = _GEN_3307 == 10'h268 ? 1'h0 : _GEN_3307 == 10'h267 | _GEN_1324; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1328 = _GEN_3307 == 10'h269 ? 1'h0 : _GEN_3307 == 10'h268 | _GEN_1326; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1330 = _GEN_3307 == 10'h26a ? 1'h0 : _GEN_3307 == 10'h269 | _GEN_1328; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1332 = _GEN_3307 == 10'h26b ? 1'h0 : _GEN_3307 == 10'h26a | _GEN_1330; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1334 = _GEN_3307 == 10'h26c ? 1'h0 : _GEN_3307 == 10'h26b | _GEN_1332; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1336 = _GEN_3307 == 10'h26d ? 1'h0 : _GEN_3307 == 10'h26c | _GEN_1334; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1338 = _GEN_3307 == 10'h26e ? 1'h0 : _GEN_3307 == 10'h26d | _GEN_1336; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1340 = _GEN_3307 == 10'h26f ? 1'h0 : _GEN_3307 == 10'h26e | _GEN_1338; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1342 = _GEN_3307 == 10'h270 ? 1'h0 : _GEN_3307 == 10'h26f | _GEN_1340; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1344 = _GEN_3307 == 10'h271 ? 1'h0 : _GEN_3307 == 10'h270 | _GEN_1342; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1346 = _GEN_3307 == 10'h272 ? 1'h0 : _GEN_3307 == 10'h271 | _GEN_1344; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1348 = _GEN_3307 == 10'h273 ? 1'h0 : _GEN_3307 == 10'h272 | _GEN_1346; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1350 = _GEN_3307 == 10'h274 ? 1'h0 : _GEN_3307 == 10'h273 | _GEN_1348; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1352 = _GEN_3307 == 10'h275 ? 1'h0 : _GEN_3307 == 10'h274 | _GEN_1350; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1354 = _GEN_3307 == 10'h276 ? 1'h0 : _GEN_3307 == 10'h275 | _GEN_1352; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1356 = _GEN_3307 == 10'h277 ? 1'h0 : _GEN_3307 == 10'h276 | _GEN_1354; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1358 = _GEN_3307 == 10'h278 ? 1'h0 : _GEN_3307 == 10'h277 | _GEN_1356; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1360 = _GEN_3307 == 10'h279 ? 1'h0 : _GEN_3307 == 10'h278 | _GEN_1358; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1362 = _GEN_3307 == 10'h27a ? 1'h0 : _GEN_3307 == 10'h279 | _GEN_1360; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1364 = _GEN_3307 == 10'h27b ? 1'h0 : _GEN_3307 == 10'h27a | _GEN_1362; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1366 = _GEN_3307 == 10'h27c ? 1'h0 : _GEN_3307 == 10'h27b | _GEN_1364; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1368 = _GEN_3307 == 10'h27d ? 1'h0 : _GEN_3307 == 10'h27c | _GEN_1366; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1370 = _GEN_3307 == 10'h27e ? 1'h0 : _GEN_3307 == 10'h27d | _GEN_1368; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1372 = _GEN_3307 == 10'h27f ? 1'h0 : _GEN_3307 == 10'h27e | _GEN_1370; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1374 = _GEN_3307 == 10'h280 ? 1'h0 : _GEN_3307 == 10'h27f | _GEN_1372; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1376 = _GEN_3307 == 10'h281 ? 1'h0 : _GEN_3307 == 10'h280 | _GEN_1374; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1378 = _GEN_3307 == 10'h282 ? 1'h0 : _GEN_3307 == 10'h281 | _GEN_1376; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1380 = _GEN_3307 == 10'h283 ? 1'h0 : _GEN_3307 == 10'h282 | _GEN_1378; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1382 = _GEN_3307 == 10'h284 ? 1'h0 : _GEN_3307 == 10'h283 | _GEN_1380; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1384 = _GEN_3307 == 10'h285 ? 1'h0 : _GEN_3307 == 10'h284 | _GEN_1382; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1386 = _GEN_3307 == 10'h286 ? 1'h0 : _GEN_3307 == 10'h285 | _GEN_1384; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1388 = _GEN_3307 == 10'h287 ? 1'h0 : _GEN_3307 == 10'h286 | _GEN_1386; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1390 = _GEN_3307 == 10'h288 ? 1'h0 : _GEN_3307 == 10'h287 | _GEN_1388; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1392 = _GEN_3307 == 10'h289 ? 1'h0 : _GEN_3307 == 10'h288 | _GEN_1390; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1394 = _GEN_3307 == 10'h28a ? 1'h0 : _GEN_3307 == 10'h289 | _GEN_1392; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1396 = _GEN_3307 == 10'h28b ? 1'h0 : _GEN_3307 == 10'h28a | _GEN_1394; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1398 = _GEN_3307 == 10'h28c ? 1'h0 : _GEN_3307 == 10'h28b | _GEN_1396; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1400 = _GEN_3307 == 10'h28d ? 1'h0 : _GEN_3307 == 10'h28c | _GEN_1398; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1402 = _GEN_3307 == 10'h28e ? 1'h0 : _GEN_3307 == 10'h28d | _GEN_1400; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1404 = _GEN_3307 == 10'h28f ? 1'h0 : _GEN_3307 == 10'h28e | _GEN_1402; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1406 = _GEN_3307 == 10'h290 ? 1'h0 : _GEN_3307 == 10'h28f | _GEN_1404; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1408 = _GEN_3307 == 10'h291 ? 1'h0 : _GEN_3307 == 10'h290 | _GEN_1406; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1410 = _GEN_3307 == 10'h292 ? 1'h0 : _GEN_3307 == 10'h291 | _GEN_1408; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1412 = _GEN_3307 == 10'h293 ? 1'h0 : _GEN_3307 == 10'h292 | _GEN_1410; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1414 = _GEN_3307 == 10'h294 ? 1'h0 : _GEN_3307 == 10'h293 | _GEN_1412; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1416 = i == 8'h0 ? 1'h0 : _GEN_1158; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1417 = i == 8'h1 ? 1'h0 : _GEN_1416; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1418 = i == 8'h4 ? 1'h0 : _GEN_1417; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1421 = i == 8'h2b ? 1'h0 : i == 8'h16 | (i == 8'h15 | _GEN_1418); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1422 = i == 8'h2e ? 1'h0 : _GEN_1421; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1423 = i == 8'h58 ? 1'h0 : _GEN_1422; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1424 = i == 8'h5d ? 1'h0 : _GEN_1423; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1425 = i == 8'hb2 ? 1'h0 : _GEN_1424; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1427 = _GEN_3306 == 9'h166 ? 1'h0 : i == 8'hbb | _GEN_1425; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1431 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_3307 == 10'h2f2 | (_GEN_3306 == 9'h178 | (_GEN_3306 == 9'h166 |
    _GEN_1427)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1432 = i == 8'h1 ? 1'h0 : _GEN_1176; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1433 = i == 8'h2 ? 1'h0 : _GEN_1432; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1434 = i == 8'h5 ? 1'h0 : _GEN_1433; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1435 = i == 8'h9 ? 1'h0 : _GEN_1434; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1436 = i == 8'hb ? 1'h0 : _GEN_1435; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1437 = i == 8'h14 ? 1'h0 : _GEN_1436; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1438 = i == 8'h17 ? 1'h0 : _GEN_1437; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1439 = i == 8'h2a ? 1'h0 : _GEN_1438; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1441 = i == 8'h2c ? 1'h0 : i == 8'h2b | _GEN_1439; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1442 = i == 8'h2d ? 1'h0 : _GEN_1441; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1444 = i == 8'h2f ? 1'h0 : i == 8'h2e | _GEN_1442; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1445 = i == 8'h56 ? 1'h0 : _GEN_1444; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1447 = i == 8'h5a ? 1'h0 : i == 8'h58 | _GEN_1445; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1448 = i == 8'h5b ? 1'h0 : _GEN_1447; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1450 = i == 8'h5f ? 1'h0 : i == 8'h5d | _GEN_1448; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1451 = i == 8'hae ? 1'h0 : _GEN_1450; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1453 = i == 8'hb6 ? 1'h0 : i == 8'hb2 | _GEN_1451; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1455 = i == 8'hbb ? 1'h0 : i == 8'hb7 | _GEN_1453; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1457 = _GEN_3306 == 9'h15e ? 1'h0 : i == 8'hbf | _GEN_1455; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1460 = _GEN_3306 == 9'h166 ? 1'h0 : _GEN_3306 == 9'h166 | (_GEN_3306 == 9'h15e | _GEN_1457); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1461 = _GEN_3306 == 9'h16e ? 1'h0 : _GEN_1460; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1464 = _GEN_3306 == 9'h178 ? 1'h0 : _GEN_3306 == 9'h170 | (_GEN_3306 == 9'h16e | _GEN_1461); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1467 = _GEN_3307 == 10'h2e2 ? 1'h0 : _GEN_3307 == 10'h2e2 | (_GEN_3306 == 9'h180 | _GEN_1464); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1468 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_1467; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1471 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_3307 == 10'h302 | (_GEN_3307 == 10'h2f2 | _GEN_1468); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1472 = i == 8'h1 ? 1'h0 : _GEN_1195; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1473 = i == 8'h2 ? 1'h0 : _GEN_1472; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1474 = i == 8'h5 ? 1'h0 : _GEN_1473; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1475 = i == 8'h9 ? 1'h0 : _GEN_1474; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1476 = i == 8'hb ? 1'h0 : _GEN_1475; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1477 = i == 8'h14 ? 1'h0 : _GEN_1476; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1478 = i == 8'h17 ? 1'h0 : _GEN_1477; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1479 = i == 8'h55 ? 1'h0 : _GEN_1478; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1481 = i == 8'h57 ? 1'h0 : i == 8'h56 | _GEN_1479; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1483 = i == 8'h59 ? 1'h0 : i == 8'h58 | _GEN_1481; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1486 = i == 8'h5c ? 1'h0 : i == 8'h5b | (i == 8'h5a | _GEN_1483); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1488 = i == 8'h5e ? 1'h0 : i == 8'h5d | _GEN_1486; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1490 = i == 8'h60 ? 1'h0 : i == 8'h5f | _GEN_1488; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1491 = i == 8'hac ? 1'h0 : _GEN_1490; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1493 = i == 8'hb0 ? 1'h0 : i == 8'hae | _GEN_1491; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1495 = i == 8'hb4 ? 1'h0 : i == 8'hb2 | _GEN_1493; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1497 = i == 8'hb7 ? 1'h0 : i == 8'hb6 | _GEN_1495; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1499 = i == 8'hbb ? 1'h0 : i == 8'hb9 | _GEN_1497; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1501 = i == 8'hbf ? 1'h0 : i == 8'hbd | _GEN_1499; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1503 = _GEN_3306 == 9'h15a ? 1'h0 : i == 8'hc1 | _GEN_1501; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1506 = _GEN_3306 == 9'h15e ? 1'h0 : _GEN_3306 == 9'h15e | (_GEN_3306 == 9'h15a | _GEN_1503); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1507 = _GEN_3306 == 9'h162 ? 1'h0 : _GEN_1506; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1510 = _GEN_3306 == 9'h166 ? 1'h0 : _GEN_3306 == 9'h166 | (_GEN_3306 == 9'h162 | _GEN_1507); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1511 = _GEN_3306 == 9'h16a ? 1'h0 : _GEN_1510; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1514 = _GEN_3306 == 9'h16e ? 1'h0 : _GEN_3306 == 9'h16e | (_GEN_3306 == 9'h16a | _GEN_1511); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1515 = _GEN_3306 == 9'h170 ? 1'h0 : _GEN_1514; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1517 = _GEN_3306 == 9'h178 ? 1'h0 : _GEN_3306 == 9'h174 | _GEN_1515; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1519 = _GEN_3306 == 9'h180 ? 1'h0 : _GEN_3306 == 9'h17c | _GEN_1517; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1521 = _GEN_3307 == 10'h2e2 ? 1'h0 : _GEN_3306 == 9'h184 | _GEN_1519; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1524 = _GEN_3307 == 10'h2ea ? 1'h0 : _GEN_3307 == 10'h2ea | (_GEN_3307 == 10'h2e2 | _GEN_1521); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1525 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_1524; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1528 = _GEN_3307 == 10'h2fa ? 1'h0 : _GEN_3307 == 10'h2fa | (_GEN_3307 == 10'h2f2 | _GEN_1525); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1529 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_1528; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1532 = _GEN_3307 == 10'h30a ? 1'h0 : _GEN_3307 == 10'h30a | (_GEN_3307 == 10'h302 | _GEN_1529); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1533 = i == 8'h1 ? 1'h0 : _GEN_1214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1534 = i == 8'h2 ? 1'h0 : _GEN_1533; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1535 = i == 8'h5 ? 1'h0 : _GEN_1534; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1536 = i == 8'h9 ? 1'h0 : _GEN_1535; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1537 = i == 8'hb ? 1'h0 : _GEN_1536; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1538 = i == 8'h14 ? 1'h0 : _GEN_1537; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1539 = i == 8'h17 ? 1'h0 : _GEN_1538; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1540 = i == 8'hab ? 1'h0 : _GEN_1539; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1542 = i == 8'had ? 1'h0 : i == 8'hac | _GEN_1540; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1544 = i == 8'haf ? 1'h0 : i == 8'hae | _GEN_1542; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1546 = i == 8'hb1 ? 1'h0 : i == 8'hb0 | _GEN_1544; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1548 = i == 8'hb3 ? 1'h0 : i == 8'hb2 | _GEN_1546; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1550 = i == 8'hb5 ? 1'h0 : i == 8'hb4 | _GEN_1548; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1552 = i == 8'hb7 ? 1'h0 : i == 8'hb6 | _GEN_1550; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1554 = i == 8'hb9 ? 1'h0 : i == 8'hb8 | _GEN_1552; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1556 = i == 8'hbb ? 1'h0 : i == 8'hba | _GEN_1554; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1558 = i == 8'hbd ? 1'h0 : i == 8'hbc | _GEN_1556; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1560 = i == 8'hbf ? 1'h0 : i == 8'hbe | _GEN_1558; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1562 = i == 8'hc1 ? 1'h0 : i == 8'hc0 | _GEN_1560; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1564 = _GEN_3306 == 9'h158 ? 1'h0 : i == 8'hc2 | _GEN_1562; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1567 = _GEN_3306 == 9'h15a ? 1'h0 : _GEN_3306 == 9'h15a | (_GEN_3306 == 9'h158 | _GEN_1564); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1568 = _GEN_3306 == 9'h15c ? 1'h0 : _GEN_1567; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1571 = _GEN_3306 == 9'h15e ? 1'h0 : _GEN_3306 == 9'h15e | (_GEN_3306 == 9'h15c | _GEN_1568); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1572 = _GEN_3306 == 9'h160 ? 1'h0 : _GEN_1571; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1575 = _GEN_3306 == 9'h162 ? 1'h0 : _GEN_3306 == 9'h162 | (_GEN_3306 == 9'h160 | _GEN_1572); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1576 = _GEN_3306 == 9'h164 ? 1'h0 : _GEN_1575; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1579 = _GEN_3306 == 9'h166 ? 1'h0 : _GEN_3306 == 9'h166 | (_GEN_3306 == 9'h164 | _GEN_1576); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1580 = _GEN_3306 == 9'h168 ? 1'h0 : _GEN_1579; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1583 = _GEN_3306 == 9'h16a ? 1'h0 : _GEN_3306 == 9'h16a | (_GEN_3306 == 9'h168 | _GEN_1580); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1584 = _GEN_3306 == 9'h16c ? 1'h0 : _GEN_1583; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1587 = _GEN_3306 == 9'h16e ? 1'h0 : _GEN_3306 == 9'h16e | (_GEN_3306 == 9'h16c | _GEN_1584); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1588 = _GEN_3306 == 9'h170 ? 1'h0 : _GEN_1587; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1590 = _GEN_3306 == 9'h174 ? 1'h0 : _GEN_3306 == 9'h172 | _GEN_1588; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1592 = _GEN_3306 == 9'h178 ? 1'h0 : _GEN_3306 == 9'h176 | _GEN_1590; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1594 = _GEN_3306 == 9'h17c ? 1'h0 : _GEN_3306 == 9'h17a | _GEN_1592; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1596 = _GEN_3306 == 9'h180 ? 1'h0 : _GEN_3306 == 9'h17e | _GEN_1594; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1598 = _GEN_3306 == 9'h184 ? 1'h0 : _GEN_3306 == 9'h182 | _GEN_1596; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1600 = _GEN_3307 == 10'h2e2 ? 1'h0 : _GEN_3306 == 9'h186 | _GEN_1598; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1603 = _GEN_3307 == 10'h2e6 ? 1'h0 : _GEN_3307 == 10'h2e6 | (_GEN_3307 == 10'h2e2 | _GEN_1600); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1604 = _GEN_3307 == 10'h2ea ? 1'h0 : _GEN_1603; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1607 = _GEN_3307 == 10'h2ee ? 1'h0 : _GEN_3307 == 10'h2ee | (_GEN_3307 == 10'h2ea | _GEN_1604); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1608 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_1607; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1611 = _GEN_3307 == 10'h2f6 ? 1'h0 : _GEN_3307 == 10'h2f6 | (_GEN_3307 == 10'h2f2 | _GEN_1608); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1612 = _GEN_3307 == 10'h2fa ? 1'h0 : _GEN_1611; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1615 = _GEN_3307 == 10'h2fe ? 1'h0 : _GEN_3307 == 10'h2fe | (_GEN_3307 == 10'h2fa | _GEN_1612); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1616 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_1615; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1619 = _GEN_3307 == 10'h306 ? 1'h0 : _GEN_3307 == 10'h306 | (_GEN_3307 == 10'h302 | _GEN_1616); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1620 = _GEN_3307 == 10'h30a ? 1'h0 : _GEN_1619; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1623 = _GEN_3307 == 10'h30e ? 1'h0 : _GEN_3307 == 10'h30e | (_GEN_3307 == 10'h30a | _GEN_1620); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1624 = i == 8'h1 ? 1'h0 : _GEN_1249; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1625 = i == 8'h2 ? 1'h0 : _GEN_1624; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1626 = i == 8'h5 ? 1'h0 : _GEN_1625; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1627 = i == 8'h9 ? 1'h0 : _GEN_1626; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1628 = i == 8'hb ? 1'h0 : _GEN_1627; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1629 = i == 8'h14 ? 1'h0 : _GEN_1628; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1630 = i == 8'h30 ? 1'h0 : _GEN_1629; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1631 = i == 8'h61 ? 1'h0 : _GEN_1630; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1632 = i == 8'hc3 ? 1'h0 : _GEN_1631; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1633 = _GEN_3306 == 9'h157 ? 1'h0 : _GEN_1632; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1636 = _GEN_3306 == 9'h158 ? 1'h0 : _GEN_3306 == 9'h158 | (_GEN_3306 == 9'h157 | _GEN_1633); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1637 = _GEN_3306 == 9'h159 ? 1'h0 : _GEN_1636; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1640 = _GEN_3306 == 9'h15a ? 1'h0 : _GEN_3306 == 9'h15a | (_GEN_3306 == 9'h159 | _GEN_1637); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1641 = _GEN_3306 == 9'h15b ? 1'h0 : _GEN_1640; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1644 = _GEN_3306 == 9'h15c ? 1'h0 : _GEN_3306 == 9'h15c | (_GEN_3306 == 9'h15b | _GEN_1641); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1645 = _GEN_3306 == 9'h15d ? 1'h0 : _GEN_1644; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1648 = _GEN_3306 == 9'h15e ? 1'h0 : _GEN_3306 == 9'h15e | (_GEN_3306 == 9'h15d | _GEN_1645); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1649 = _GEN_3306 == 9'h15f ? 1'h0 : _GEN_1648; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1652 = _GEN_3306 == 9'h160 ? 1'h0 : _GEN_3306 == 9'h160 | (_GEN_3306 == 9'h15f | _GEN_1649); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1653 = _GEN_3306 == 9'h161 ? 1'h0 : _GEN_1652; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1656 = _GEN_3306 == 9'h162 ? 1'h0 : _GEN_3306 == 9'h162 | (_GEN_3306 == 9'h161 | _GEN_1653); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1657 = _GEN_3306 == 9'h163 ? 1'h0 : _GEN_1656; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1660 = _GEN_3306 == 9'h164 ? 1'h0 : _GEN_3306 == 9'h164 | (_GEN_3306 == 9'h163 | _GEN_1657); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1661 = _GEN_3306 == 9'h165 ? 1'h0 : _GEN_1660; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1664 = _GEN_3306 == 9'h166 ? 1'h0 : _GEN_3306 == 9'h166 | (_GEN_3306 == 9'h165 | _GEN_1661); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1665 = _GEN_3306 == 9'h167 ? 1'h0 : _GEN_1664; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1668 = _GEN_3306 == 9'h168 ? 1'h0 : _GEN_3306 == 9'h168 | (_GEN_3306 == 9'h167 | _GEN_1665); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1669 = _GEN_3306 == 9'h169 ? 1'h0 : _GEN_1668; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1672 = _GEN_3306 == 9'h16a ? 1'h0 : _GEN_3306 == 9'h16a | (_GEN_3306 == 9'h169 | _GEN_1669); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1673 = _GEN_3306 == 9'h16b ? 1'h0 : _GEN_1672; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1676 = _GEN_3306 == 9'h16c ? 1'h0 : _GEN_3306 == 9'h16c | (_GEN_3306 == 9'h16b | _GEN_1673); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1677 = _GEN_3306 == 9'h16d ? 1'h0 : _GEN_1676; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1680 = _GEN_3306 == 9'h16e ? 1'h0 : _GEN_3306 == 9'h16e | (_GEN_3306 == 9'h16d | _GEN_1677); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1681 = _GEN_3306 == 9'h16f ? 1'h0 : _GEN_1680; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1682 = _GEN_3306 == 9'h170 ? 1'h0 : _GEN_1681; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1684 = _GEN_3306 == 9'h172 ? 1'h0 : _GEN_3306 == 9'h171 | _GEN_1682; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1686 = _GEN_3306 == 9'h174 ? 1'h0 : _GEN_3306 == 9'h173 | _GEN_1684; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1688 = _GEN_3306 == 9'h176 ? 1'h0 : _GEN_3306 == 9'h175 | _GEN_1686; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1690 = _GEN_3306 == 9'h178 ? 1'h0 : _GEN_3306 == 9'h177 | _GEN_1688; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1692 = _GEN_3306 == 9'h17a ? 1'h0 : _GEN_3306 == 9'h179 | _GEN_1690; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1694 = _GEN_3306 == 9'h17c ? 1'h0 : _GEN_3306 == 9'h17b | _GEN_1692; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1696 = _GEN_3306 == 9'h17e ? 1'h0 : _GEN_3306 == 9'h17d | _GEN_1694; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1698 = _GEN_3306 == 9'h180 ? 1'h0 : _GEN_3306 == 9'h17f | _GEN_1696; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1700 = _GEN_3306 == 9'h182 ? 1'h0 : _GEN_3306 == 9'h181 | _GEN_1698; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1702 = _GEN_3306 == 9'h184 ? 1'h0 : _GEN_3306 == 9'h183 | _GEN_1700; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1704 = _GEN_3306 == 9'h186 ? 1'h0 : _GEN_3306 == 9'h185 | _GEN_1702; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1707 = _GEN_3307 == 10'h2e0 ? 1'h0 : _GEN_3307 == 10'h2e0 | (_GEN_3306 == 9'h187 | _GEN_1704); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1708 = _GEN_3307 == 10'h2e2 ? 1'h0 : _GEN_1707; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1711 = _GEN_3307 == 10'h2e4 ? 1'h0 : _GEN_3307 == 10'h2e4 | (_GEN_3307 == 10'h2e2 | _GEN_1708); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1712 = _GEN_3307 == 10'h2e6 ? 1'h0 : _GEN_1711; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1715 = _GEN_3307 == 10'h2e8 ? 1'h0 : _GEN_3307 == 10'h2e8 | (_GEN_3307 == 10'h2e6 | _GEN_1712); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1716 = _GEN_3307 == 10'h2ea ? 1'h0 : _GEN_1715; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1719 = _GEN_3307 == 10'h2ec ? 1'h0 : _GEN_3307 == 10'h2ec | (_GEN_3307 == 10'h2ea | _GEN_1716); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1720 = _GEN_3307 == 10'h2ee ? 1'h0 : _GEN_1719; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1723 = _GEN_3307 == 10'h2f0 ? 1'h0 : _GEN_3307 == 10'h2f0 | (_GEN_3307 == 10'h2ee | _GEN_1720); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1724 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_1723; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1727 = _GEN_3307 == 10'h2f4 ? 1'h0 : _GEN_3307 == 10'h2f4 | (_GEN_3307 == 10'h2f2 | _GEN_1724); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1728 = _GEN_3307 == 10'h2f6 ? 1'h0 : _GEN_1727; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1731 = _GEN_3307 == 10'h2f8 ? 1'h0 : _GEN_3307 == 10'h2f8 | (_GEN_3307 == 10'h2f6 | _GEN_1728); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1732 = _GEN_3307 == 10'h2fa ? 1'h0 : _GEN_1731; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1735 = _GEN_3307 == 10'h2fc ? 1'h0 : _GEN_3307 == 10'h2fc | (_GEN_3307 == 10'h2fa | _GEN_1732); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1736 = _GEN_3307 == 10'h2fe ? 1'h0 : _GEN_1735; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1739 = _GEN_3307 == 10'h300 ? 1'h0 : _GEN_3307 == 10'h300 | (_GEN_3307 == 10'h2fe | _GEN_1736); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1740 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_1739; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1743 = _GEN_3307 == 10'h304 ? 1'h0 : _GEN_3307 == 10'h304 | (_GEN_3307 == 10'h302 | _GEN_1740); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1744 = _GEN_3307 == 10'h306 ? 1'h0 : _GEN_1743; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1747 = _GEN_3307 == 10'h308 ? 1'h0 : _GEN_3307 == 10'h308 | (_GEN_3307 == 10'h306 | _GEN_1744); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1748 = _GEN_3307 == 10'h30a ? 1'h0 : _GEN_1747; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1751 = _GEN_3307 == 10'h30c ? 1'h0 : _GEN_3307 == 10'h30c | (_GEN_3307 == 10'h30a | _GEN_1748); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1752 = _GEN_3307 == 10'h30e ? 1'h0 : _GEN_1751; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1755 = _GEN_3307 == 10'h310 ? 1'h0 : _GEN_3307 == 10'h310 | (_GEN_3307 == 10'h30e | _GEN_1752); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1756 = i == 8'h1 ? 1'h0 : _GEN_3306 == 9'h149 | _GEN_1306; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1757 = i == 8'h2 ? 1'h0 : _GEN_1756; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1758 = i == 8'h5 ? 1'h0 : _GEN_1757; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1759 = i == 8'h9 ? 1'h0 : _GEN_1758; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1760 = i == 8'hb ? 1'h0 : _GEN_1759; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1761 = i == 8'h14 ? 1'h0 : _GEN_1760; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1762 = i == 8'h30 ? 1'h0 : _GEN_1761; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1763 = i == 8'h61 ? 1'h0 : _GEN_1762; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1765 = _GEN_3306 == 9'h157 ? 1'h0 : _GEN_3306 == 9'h157 | _GEN_1763; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1767 = _GEN_3306 == 9'h158 ? 1'h0 : _GEN_3306 == 9'h158 | _GEN_1765; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1769 = _GEN_3306 == 9'h159 ? 1'h0 : _GEN_3306 == 9'h159 | _GEN_1767; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1771 = _GEN_3306 == 9'h15a ? 1'h0 : _GEN_3306 == 9'h15a | _GEN_1769; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1773 = _GEN_3306 == 9'h15b ? 1'h0 : _GEN_3306 == 9'h15b | _GEN_1771; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1775 = _GEN_3306 == 9'h15c ? 1'h0 : _GEN_3306 == 9'h15c | _GEN_1773; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1777 = _GEN_3306 == 9'h15d ? 1'h0 : _GEN_3306 == 9'h15d | _GEN_1775; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1779 = _GEN_3306 == 9'h15e ? 1'h0 : _GEN_3306 == 9'h15e | _GEN_1777; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1781 = _GEN_3306 == 9'h15f ? 1'h0 : _GEN_3306 == 9'h15f | _GEN_1779; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1783 = _GEN_3306 == 9'h160 ? 1'h0 : _GEN_3306 == 9'h160 | _GEN_1781; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1785 = _GEN_3306 == 9'h161 ? 1'h0 : _GEN_3306 == 9'h161 | _GEN_1783; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1787 = _GEN_3306 == 9'h162 ? 1'h0 : _GEN_3306 == 9'h162 | _GEN_1785; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1789 = _GEN_3306 == 9'h163 ? 1'h0 : _GEN_3306 == 9'h163 | _GEN_1787; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1791 = _GEN_3306 == 9'h164 ? 1'h0 : _GEN_3306 == 9'h164 | _GEN_1789; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1793 = _GEN_3306 == 9'h165 ? 1'h0 : _GEN_3306 == 9'h165 | _GEN_1791; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1795 = _GEN_3306 == 9'h166 ? 1'h0 : _GEN_3306 == 9'h166 | _GEN_1793; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1797 = _GEN_3306 == 9'h167 ? 1'h0 : _GEN_3306 == 9'h167 | _GEN_1795; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1799 = _GEN_3306 == 9'h168 ? 1'h0 : _GEN_3306 == 9'h168 | _GEN_1797; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1801 = _GEN_3306 == 9'h169 ? 1'h0 : _GEN_3306 == 9'h169 | _GEN_1799; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1803 = _GEN_3306 == 9'h16a ? 1'h0 : _GEN_3306 == 9'h16a | _GEN_1801; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1805 = _GEN_3306 == 9'h16b ? 1'h0 : _GEN_3306 == 9'h16b | _GEN_1803; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1807 = _GEN_3306 == 9'h16c ? 1'h0 : _GEN_3306 == 9'h16c | _GEN_1805; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1809 = _GEN_3306 == 9'h16d ? 1'h0 : _GEN_3306 == 9'h16d | _GEN_1807; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1811 = _GEN_3306 == 9'h16e ? 1'h0 : _GEN_3306 == 9'h16e | _GEN_1809; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1813 = _GEN_3306 == 9'h188 ? 1'h0 : _GEN_3306 == 9'h16f | _GEN_1811; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1814 = _GEN_3307 == 10'h2e0 ? 1'h0 : _GEN_1813; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1817 = _GEN_3307 == 10'h2e1 ? 1'h0 : _GEN_3307 == 10'h2e1 | (_GEN_3307 == 10'h2e0 | _GEN_1814); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1818 = _GEN_3307 == 10'h2e2 ? 1'h0 : _GEN_1817; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1821 = _GEN_3307 == 10'h2e3 ? 1'h0 : _GEN_3307 == 10'h2e3 | (_GEN_3307 == 10'h2e2 | _GEN_1818); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1822 = _GEN_3307 == 10'h2e4 ? 1'h0 : _GEN_1821; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1825 = _GEN_3307 == 10'h2e5 ? 1'h0 : _GEN_3307 == 10'h2e5 | (_GEN_3307 == 10'h2e4 | _GEN_1822); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1826 = _GEN_3307 == 10'h2e6 ? 1'h0 : _GEN_1825; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1829 = _GEN_3307 == 10'h2e7 ? 1'h0 : _GEN_3307 == 10'h2e7 | (_GEN_3307 == 10'h2e6 | _GEN_1826); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1830 = _GEN_3307 == 10'h2e8 ? 1'h0 : _GEN_1829; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1833 = _GEN_3307 == 10'h2e9 ? 1'h0 : _GEN_3307 == 10'h2e9 | (_GEN_3307 == 10'h2e8 | _GEN_1830); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1834 = _GEN_3307 == 10'h2ea ? 1'h0 : _GEN_1833; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1837 = _GEN_3307 == 10'h2eb ? 1'h0 : _GEN_3307 == 10'h2eb | (_GEN_3307 == 10'h2ea | _GEN_1834); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1838 = _GEN_3307 == 10'h2ec ? 1'h0 : _GEN_1837; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1841 = _GEN_3307 == 10'h2ed ? 1'h0 : _GEN_3307 == 10'h2ed | (_GEN_3307 == 10'h2ec | _GEN_1838); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1842 = _GEN_3307 == 10'h2ee ? 1'h0 : _GEN_1841; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1845 = _GEN_3307 == 10'h2ef ? 1'h0 : _GEN_3307 == 10'h2ef | (_GEN_3307 == 10'h2ee | _GEN_1842); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1846 = _GEN_3307 == 10'h2f0 ? 1'h0 : _GEN_1845; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1849 = _GEN_3307 == 10'h2f1 ? 1'h0 : _GEN_3307 == 10'h2f1 | (_GEN_3307 == 10'h2f0 | _GEN_1846); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1850 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_1849; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1853 = _GEN_3307 == 10'h2f3 ? 1'h0 : _GEN_3307 == 10'h2f3 | (_GEN_3307 == 10'h2f2 | _GEN_1850); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1854 = _GEN_3307 == 10'h2f4 ? 1'h0 : _GEN_1853; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1857 = _GEN_3307 == 10'h2f5 ? 1'h0 : _GEN_3307 == 10'h2f5 | (_GEN_3307 == 10'h2f4 | _GEN_1854); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1858 = _GEN_3307 == 10'h2f6 ? 1'h0 : _GEN_1857; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1861 = _GEN_3307 == 10'h2f7 ? 1'h0 : _GEN_3307 == 10'h2f7 | (_GEN_3307 == 10'h2f6 | _GEN_1858); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1862 = _GEN_3307 == 10'h2f8 ? 1'h0 : _GEN_1861; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1865 = _GEN_3307 == 10'h2f9 ? 1'h0 : _GEN_3307 == 10'h2f9 | (_GEN_3307 == 10'h2f8 | _GEN_1862); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1866 = _GEN_3307 == 10'h2fa ? 1'h0 : _GEN_1865; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1869 = _GEN_3307 == 10'h2fb ? 1'h0 : _GEN_3307 == 10'h2fb | (_GEN_3307 == 10'h2fa | _GEN_1866); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1870 = _GEN_3307 == 10'h2fc ? 1'h0 : _GEN_1869; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1873 = _GEN_3307 == 10'h2fd ? 1'h0 : _GEN_3307 == 10'h2fd | (_GEN_3307 == 10'h2fc | _GEN_1870); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1874 = _GEN_3307 == 10'h2fe ? 1'h0 : _GEN_1873; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1877 = _GEN_3307 == 10'h2ff ? 1'h0 : _GEN_3307 == 10'h2ff | (_GEN_3307 == 10'h2fe | _GEN_1874); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1878 = _GEN_3307 == 10'h300 ? 1'h0 : _GEN_1877; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1881 = _GEN_3307 == 10'h301 ? 1'h0 : _GEN_3307 == 10'h301 | (_GEN_3307 == 10'h300 | _GEN_1878); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1882 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_1881; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1885 = _GEN_3307 == 10'h303 ? 1'h0 : _GEN_3307 == 10'h303 | (_GEN_3307 == 10'h302 | _GEN_1882); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1886 = _GEN_3307 == 10'h304 ? 1'h0 : _GEN_1885; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1889 = _GEN_3307 == 10'h305 ? 1'h0 : _GEN_3307 == 10'h305 | (_GEN_3307 == 10'h304 | _GEN_1886); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1890 = _GEN_3307 == 10'h306 ? 1'h0 : _GEN_1889; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1893 = _GEN_3307 == 10'h307 ? 1'h0 : _GEN_3307 == 10'h307 | (_GEN_3307 == 10'h306 | _GEN_1890); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1894 = _GEN_3307 == 10'h308 ? 1'h0 : _GEN_1893; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1897 = _GEN_3307 == 10'h309 ? 1'h0 : _GEN_3307 == 10'h309 | (_GEN_3307 == 10'h308 | _GEN_1894); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1898 = _GEN_3307 == 10'h30a ? 1'h0 : _GEN_1897; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1901 = _GEN_3307 == 10'h30b ? 1'h0 : _GEN_3307 == 10'h30b | (_GEN_3307 == 10'h30a | _GEN_1898); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1902 = _GEN_3307 == 10'h30c ? 1'h0 : _GEN_1901; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1905 = _GEN_3307 == 10'h30d ? 1'h0 : _GEN_3307 == 10'h30d | (_GEN_3307 == 10'h30c | _GEN_1902); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1906 = _GEN_3307 == 10'h30e ? 1'h0 : _GEN_1905; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1909 = _GEN_3307 == 10'h30f ? 1'h0 : _GEN_3307 == 10'h30f | (_GEN_3307 == 10'h30e | _GEN_1906); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1910 = _GEN_3307 == 10'h310 ? 1'h0 : _GEN_1909; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1913 = _GEN_3307 == 10'h311 ? 1'h0 : _GEN_3307 == 10'h311 | (_GEN_3307 == 10'h310 | _GEN_1910); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1914 = i == 8'h1 ? 1'h0 : _GEN_3307 == 10'h294 | _GEN_1414; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1915 = i == 8'h2 ? 1'h0 : _GEN_1914; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1916 = i == 8'h5 ? 1'h0 : _GEN_1915; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1917 = i == 8'h9 ? 1'h0 : _GEN_1916; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1918 = i == 8'hb ? 1'h0 : _GEN_1917; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1919 = i == 8'h29 ? 1'h0 : _GEN_1918; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1920 = i == 8'h30 ? 1'h0 : _GEN_1919; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1921 = i == 8'h54 ? 1'h0 : _GEN_1920; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1922 = i == 8'h61 ? 1'h0 : _GEN_1921; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1923 = i == 8'haa ? 1'h0 : _GEN_1922; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1924 = _GEN_3306 == 9'h156 ? 1'h0 : _GEN_1923; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1925 = _GEN_3306 == 9'h188 ? 1'h0 : _GEN_1924; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1926 = _GEN_3307 == 10'h2ae ? 1'h0 : _GEN_1925; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1928 = _GEN_3307 == 10'h2af ? 1'h0 : _GEN_3307 == 10'h2ae | _GEN_1926; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1930 = _GEN_3307 == 10'h2b0 ? 1'h0 : _GEN_3307 == 10'h2af | _GEN_1928; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1932 = _GEN_3307 == 10'h2b1 ? 1'h0 : _GEN_3307 == 10'h2b0 | _GEN_1930; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1934 = _GEN_3307 == 10'h2b2 ? 1'h0 : _GEN_3307 == 10'h2b1 | _GEN_1932; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1936 = _GEN_3307 == 10'h2b3 ? 1'h0 : _GEN_3307 == 10'h2b2 | _GEN_1934; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1938 = _GEN_3307 == 10'h2b4 ? 1'h0 : _GEN_3307 == 10'h2b3 | _GEN_1936; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1940 = _GEN_3307 == 10'h2b5 ? 1'h0 : _GEN_3307 == 10'h2b4 | _GEN_1938; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1942 = _GEN_3307 == 10'h2b6 ? 1'h0 : _GEN_3307 == 10'h2b5 | _GEN_1940; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1944 = _GEN_3307 == 10'h2b7 ? 1'h0 : _GEN_3307 == 10'h2b6 | _GEN_1942; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1946 = _GEN_3307 == 10'h2b8 ? 1'h0 : _GEN_3307 == 10'h2b7 | _GEN_1944; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1948 = _GEN_3307 == 10'h2b9 ? 1'h0 : _GEN_3307 == 10'h2b8 | _GEN_1946; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1950 = _GEN_3307 == 10'h2ba ? 1'h0 : _GEN_3307 == 10'h2b9 | _GEN_1948; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1952 = _GEN_3307 == 10'h2bb ? 1'h0 : _GEN_3307 == 10'h2ba | _GEN_1950; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1954 = _GEN_3307 == 10'h2bc ? 1'h0 : _GEN_3307 == 10'h2bb | _GEN_1952; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1956 = _GEN_3307 == 10'h2bd ? 1'h0 : _GEN_3307 == 10'h2bc | _GEN_1954; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1958 = _GEN_3307 == 10'h2be ? 1'h0 : _GEN_3307 == 10'h2bd | _GEN_1956; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1960 = _GEN_3307 == 10'h2bf ? 1'h0 : _GEN_3307 == 10'h2be | _GEN_1958; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1962 = _GEN_3307 == 10'h2c0 ? 1'h0 : _GEN_3307 == 10'h2bf | _GEN_1960; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1964 = _GEN_3307 == 10'h2c1 ? 1'h0 : _GEN_3307 == 10'h2c0 | _GEN_1962; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1966 = _GEN_3307 == 10'h2c2 ? 1'h0 : _GEN_3307 == 10'h2c1 | _GEN_1964; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1968 = _GEN_3307 == 10'h2c3 ? 1'h0 : _GEN_3307 == 10'h2c2 | _GEN_1966; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1970 = _GEN_3307 == 10'h2c4 ? 1'h0 : _GEN_3307 == 10'h2c3 | _GEN_1968; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1972 = _GEN_3307 == 10'h2c5 ? 1'h0 : _GEN_3307 == 10'h2c4 | _GEN_1970; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1974 = _GEN_3307 == 10'h2c6 ? 1'h0 : _GEN_3307 == 10'h2c5 | _GEN_1972; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1976 = _GEN_3307 == 10'h2c7 ? 1'h0 : _GEN_3307 == 10'h2c6 | _GEN_1974; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1978 = _GEN_3307 == 10'h2c8 ? 1'h0 : _GEN_3307 == 10'h2c7 | _GEN_1976; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1980 = _GEN_3307 == 10'h2c9 ? 1'h0 : _GEN_3307 == 10'h2c8 | _GEN_1978; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1982 = _GEN_3307 == 10'h2ca ? 1'h0 : _GEN_3307 == 10'h2c9 | _GEN_1980; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1984 = _GEN_3307 == 10'h2cb ? 1'h0 : _GEN_3307 == 10'h2ca | _GEN_1982; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1986 = _GEN_3307 == 10'h2cc ? 1'h0 : _GEN_3307 == 10'h2cb | _GEN_1984; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1988 = _GEN_3307 == 10'h2cd ? 1'h0 : _GEN_3307 == 10'h2cc | _GEN_1986; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1990 = _GEN_3307 == 10'h2ce ? 1'h0 : _GEN_3307 == 10'h2cd | _GEN_1988; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1992 = _GEN_3307 == 10'h2cf ? 1'h0 : _GEN_3307 == 10'h2ce | _GEN_1990; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1994 = _GEN_3307 == 10'h2d0 ? 1'h0 : _GEN_3307 == 10'h2cf | _GEN_1992; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1996 = _GEN_3307 == 10'h2d1 ? 1'h0 : _GEN_3307 == 10'h2d0 | _GEN_1994; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_1998 = _GEN_3307 == 10'h2d2 ? 1'h0 : _GEN_3307 == 10'h2d1 | _GEN_1996; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2000 = _GEN_3307 == 10'h2d3 ? 1'h0 : _GEN_3307 == 10'h2d2 | _GEN_1998; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2002 = _GEN_3307 == 10'h2d4 ? 1'h0 : _GEN_3307 == 10'h2d3 | _GEN_2000; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2004 = _GEN_3307 == 10'h2d5 ? 1'h0 : _GEN_3307 == 10'h2d4 | _GEN_2002; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2006 = _GEN_3307 == 10'h2d6 ? 1'h0 : _GEN_3307 == 10'h2d5 | _GEN_2004; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2008 = _GEN_3307 == 10'h2d7 ? 1'h0 : _GEN_3307 == 10'h2d6 | _GEN_2006; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2010 = _GEN_3307 == 10'h2d8 ? 1'h0 : _GEN_3307 == 10'h2d7 | _GEN_2008; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2012 = _GEN_3307 == 10'h2d9 ? 1'h0 : _GEN_3307 == 10'h2d8 | _GEN_2010; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2014 = _GEN_3307 == 10'h2da ? 1'h0 : _GEN_3307 == 10'h2d9 | _GEN_2012; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2016 = _GEN_3307 == 10'h2db ? 1'h0 : _GEN_3307 == 10'h2da | _GEN_2014; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2018 = _GEN_3307 == 10'h2dc ? 1'h0 : _GEN_3307 == 10'h2db | _GEN_2016; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2020 = _GEN_3307 == 10'h2dd ? 1'h0 : _GEN_3307 == 10'h2dc | _GEN_2018; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2022 = _GEN_3307 == 10'h2de ? 1'h0 : _GEN_3307 == 10'h2dd | _GEN_2020; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2024 = _GEN_3307 == 10'h2df ? 1'h0 : _GEN_3307 == 10'h2de | _GEN_2022; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2026 = _GEN_3307 == 10'h2e0 ? 1'h0 : _GEN_3307 == 10'h2df | _GEN_2024; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2028 = _GEN_3307 == 10'h2e1 ? 1'h0 : _GEN_3307 == 10'h2e0 | _GEN_2026; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2030 = _GEN_3307 == 10'h2e2 ? 1'h0 : _GEN_3307 == 10'h2e1 | _GEN_2028; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2032 = _GEN_3307 == 10'h2e3 ? 1'h0 : _GEN_3307 == 10'h2e2 | _GEN_2030; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2034 = _GEN_3307 == 10'h2e4 ? 1'h0 : _GEN_3307 == 10'h2e3 | _GEN_2032; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2036 = _GEN_3307 == 10'h2e5 ? 1'h0 : _GEN_3307 == 10'h2e4 | _GEN_2034; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2038 = _GEN_3307 == 10'h2e6 ? 1'h0 : _GEN_3307 == 10'h2e5 | _GEN_2036; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2040 = _GEN_3307 == 10'h2e7 ? 1'h0 : _GEN_3307 == 10'h2e6 | _GEN_2038; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2042 = _GEN_3307 == 10'h2e8 ? 1'h0 : _GEN_3307 == 10'h2e7 | _GEN_2040; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2044 = _GEN_3307 == 10'h2e9 ? 1'h0 : _GEN_3307 == 10'h2e8 | _GEN_2042; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2046 = _GEN_3307 == 10'h2ea ? 1'h0 : _GEN_3307 == 10'h2e9 | _GEN_2044; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2048 = _GEN_3307 == 10'h2eb ? 1'h0 : _GEN_3307 == 10'h2ea | _GEN_2046; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2050 = _GEN_3307 == 10'h2ec ? 1'h0 : _GEN_3307 == 10'h2eb | _GEN_2048; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2052 = _GEN_3307 == 10'h2ed ? 1'h0 : _GEN_3307 == 10'h2ec | _GEN_2050; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2054 = _GEN_3307 == 10'h2ee ? 1'h0 : _GEN_3307 == 10'h2ed | _GEN_2052; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2056 = _GEN_3307 == 10'h2ef ? 1'h0 : _GEN_3307 == 10'h2ee | _GEN_2054; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2058 = _GEN_3307 == 10'h2f0 ? 1'h0 : _GEN_3307 == 10'h2ef | _GEN_2056; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2060 = _GEN_3307 == 10'h2f1 ? 1'h0 : _GEN_3307 == 10'h2f0 | _GEN_2058; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2062 = _GEN_3307 == 10'h2f2 ? 1'h0 : _GEN_3307 == 10'h2f1 | _GEN_2060; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2064 = _GEN_3307 == 10'h2f3 ? 1'h0 : _GEN_3307 == 10'h2f2 | _GEN_2062; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2066 = _GEN_3307 == 10'h2f4 ? 1'h0 : _GEN_3307 == 10'h2f3 | _GEN_2064; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2068 = _GEN_3307 == 10'h2f5 ? 1'h0 : _GEN_3307 == 10'h2f4 | _GEN_2066; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2070 = _GEN_3307 == 10'h2f6 ? 1'h0 : _GEN_3307 == 10'h2f5 | _GEN_2068; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2072 = _GEN_3307 == 10'h2f7 ? 1'h0 : _GEN_3307 == 10'h2f6 | _GEN_2070; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2074 = _GEN_3307 == 10'h2f8 ? 1'h0 : _GEN_3307 == 10'h2f7 | _GEN_2072; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2076 = _GEN_3307 == 10'h2f9 ? 1'h0 : _GEN_3307 == 10'h2f8 | _GEN_2074; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2078 = _GEN_3307 == 10'h2fa ? 1'h0 : _GEN_3307 == 10'h2f9 | _GEN_2076; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2080 = _GEN_3307 == 10'h2fb ? 1'h0 : _GEN_3307 == 10'h2fa | _GEN_2078; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2082 = _GEN_3307 == 10'h2fc ? 1'h0 : _GEN_3307 == 10'h2fb | _GEN_2080; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2084 = _GEN_3307 == 10'h2fd ? 1'h0 : _GEN_3307 == 10'h2fc | _GEN_2082; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2086 = _GEN_3307 == 10'h2fe ? 1'h0 : _GEN_3307 == 10'h2fd | _GEN_2084; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2088 = _GEN_3307 == 10'h2ff ? 1'h0 : _GEN_3307 == 10'h2fe | _GEN_2086; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2090 = _GEN_3307 == 10'h300 ? 1'h0 : _GEN_3307 == 10'h2ff | _GEN_2088; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2092 = _GEN_3307 == 10'h301 ? 1'h0 : _GEN_3307 == 10'h300 | _GEN_2090; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2094 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_3307 == 10'h301 | _GEN_2092; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2096 = _GEN_3307 == 10'h303 ? 1'h0 : _GEN_3307 == 10'h302 | _GEN_2094; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2098 = _GEN_3307 == 10'h304 ? 1'h0 : _GEN_3307 == 10'h303 | _GEN_2096; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2100 = _GEN_3307 == 10'h305 ? 1'h0 : _GEN_3307 == 10'h304 | _GEN_2098; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2102 = _GEN_3307 == 10'h306 ? 1'h0 : _GEN_3307 == 10'h305 | _GEN_2100; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2104 = _GEN_3307 == 10'h307 ? 1'h0 : _GEN_3307 == 10'h306 | _GEN_2102; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2106 = _GEN_3307 == 10'h308 ? 1'h0 : _GEN_3307 == 10'h307 | _GEN_2104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2108 = _GEN_3307 == 10'h309 ? 1'h0 : _GEN_3307 == 10'h308 | _GEN_2106; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2110 = _GEN_3307 == 10'h30a ? 1'h0 : _GEN_3307 == 10'h309 | _GEN_2108; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2112 = _GEN_3307 == 10'h30b ? 1'h0 : _GEN_3307 == 10'h30a | _GEN_2110; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2114 = _GEN_3307 == 10'h30c ? 1'h0 : _GEN_3307 == 10'h30b | _GEN_2112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2116 = _GEN_3307 == 10'h30d ? 1'h0 : _GEN_3307 == 10'h30c | _GEN_2114; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2118 = _GEN_3307 == 10'h30e ? 1'h0 : _GEN_3307 == 10'h30d | _GEN_2116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2120 = _GEN_3307 == 10'h30f ? 1'h0 : _GEN_3307 == 10'h30e | _GEN_2118; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2122 = _GEN_3307 == 10'h310 ? 1'h0 : _GEN_3307 == 10'h30f | _GEN_2120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2124 = _GEN_3307 == 10'h311 ? 1'h0 : _GEN_3307 == 10'h310 | _GEN_2122; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2126 = i == 8'h0 ? 1'h0 : _GEN_1431; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2130 = i == 8'h17 ? 1'h0 : i == 8'hb | (i == 8'h5 | (i == 8'h2 | _GEN_2126)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2131 = i == 8'h30 ? 1'h0 : _GEN_2130; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2133 = i == 8'hc5 ? 1'h0 : i == 8'h62 | _GEN_2131; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2135 = i == 8'h0 ? 1'h0 : _GEN_1471; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2139 = i == 8'h2f ? 1'h0 : i == 8'h18 | (i == 8'h5 | (i == 8'h2 | _GEN_2135)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2141 = i == 8'h31 ? 1'h0 : i == 8'h30 | _GEN_2139; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2143 = i == 8'h62 ? 1'h0 : i == 8'h60 | _GEN_2141; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2145 = i == 8'hc1 ? 1'h0 : i == 8'h64 | _GEN_2143; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2148 = i == 8'hc5 ? 1'h0 : i == 8'hc5 | (i == 8'hc1 | _GEN_2145); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2149 = i == 8'hc9 ? 1'h0 : _GEN_2148; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2151 = i == 8'h0 ? 1'h0 : _GEN_1532; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2152 = i == 8'h2 ? 1'h0 : _GEN_2151; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2153 = i == 8'h5 ? 1'h0 : _GEN_2152; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2154 = i == 8'h18 ? 1'h0 : _GEN_2153; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2156 = i == 8'h60 ? 1'h0 : i == 8'h5f | _GEN_2154; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2158 = i == 8'h62 ? 1'h0 : i == 8'h61 | _GEN_2156; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2160 = i == 8'h64 ? 1'h0 : i == 8'h63 | _GEN_2158; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2161 = i == 8'hbf ? 1'h0 : _GEN_2160; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2164 = i == 8'hc1 ? 1'h0 : i == 8'hc1 | (i == 8'hbf | _GEN_2161); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2165 = i == 8'hc3 ? 1'h0 : _GEN_2164; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2168 = i == 8'hc5 ? 1'h0 : i == 8'hc5 | (i == 8'hc3 | _GEN_2165); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2169 = i == 8'hc7 ? 1'h0 : _GEN_2168; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2172 = i == 8'hc9 ? 1'h0 : i == 8'hc9 | (i == 8'hc7 | _GEN_2169); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2173 = i == 8'h1 ? 1'h0 : _GEN_1623; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2174 = i == 8'h2 ? 1'h0 : _GEN_2173; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2175 = i == 8'h4 ? 1'h0 : _GEN_2174; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2176 = i == 8'h5 ? 1'h0 : _GEN_2175; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2177 = i == 8'ha ? 1'h0 : _GEN_2176; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2178 = i == 8'h16 ? 1'h0 : _GEN_2177; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2179 = i == 8'h18 ? 1'h0 : _GEN_2178; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2180 = i == 8'h2e ? 1'h0 : _GEN_2179; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2181 = i == 8'h5e ? 1'h0 : _GEN_2180; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2182 = i == 8'h64 ? 1'h0 : _GEN_2181; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2183 = i == 8'hbe ? 1'h0 : _GEN_2182; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2186 = i == 8'hbf ? 1'h0 : i == 8'hbf | (i == 8'hbe | _GEN_2183); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2187 = i == 8'hc0 ? 1'h0 : _GEN_2186; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2190 = i == 8'hc1 ? 1'h0 : i == 8'hc1 | (i == 8'hc0 | _GEN_2187); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2191 = i == 8'hc2 ? 1'h0 : _GEN_2190; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2194 = i == 8'hc3 ? 1'h0 : i == 8'hc3 | (i == 8'hc2 | _GEN_2191); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2195 = i == 8'hc4 ? 1'h0 : _GEN_2194; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2198 = i == 8'hc5 ? 1'h0 : i == 8'hc5 | (i == 8'hc4 | _GEN_2195); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2199 = i == 8'hc6 ? 1'h0 : _GEN_2198; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2202 = i == 8'hc7 ? 1'h0 : i == 8'hc7 | (i == 8'hc6 | _GEN_2199); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2203 = i == 8'hc8 ? 1'h0 : _GEN_2202; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2206 = i == 8'hc9 ? 1'h0 : i == 8'hc9 | (i == 8'hc8 | _GEN_2203); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2207 = i == 8'h1 ? 1'h0 : _GEN_1755; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2209 = i == 8'h4 ? 1'h0 : i == 8'h2 | _GEN_2207; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2211 = i == 8'ha ? 1'h0 : i == 8'h5 | _GEN_2209; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2212 = i == 8'h16 ? 1'h0 : _GEN_2211; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2214 = i == 8'h2e ? 1'h0 : i == 8'h18 | _GEN_2212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2215 = i == 8'h5e ? 1'h0 : _GEN_2214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2218 = i == 8'hbe ? 1'h0 : i == 8'hbe | (i == 8'h64 | _GEN_2215); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2220 = i == 8'hbf ? 1'h0 : i == 8'hbf | _GEN_2218; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2222 = i == 8'hc0 ? 1'h0 : i == 8'hc0 | _GEN_2220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2224 = i == 8'hc1 ? 1'h0 : i == 8'hc1 | _GEN_2222; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2226 = i == 8'hc2 ? 1'h0 : i == 8'hc2 | _GEN_2224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2228 = i == 8'hc3 ? 1'h0 : i == 8'hc3 | _GEN_2226; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2230 = i == 8'hc4 ? 1'h0 : i == 8'hc4 | _GEN_2228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2232 = i == 8'hc5 ? 1'h0 : i == 8'hc5 | _GEN_2230; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2234 = i == 8'hc6 ? 1'h0 : i == 8'hc6 | _GEN_2232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2236 = i == 8'hc7 ? 1'h0 : i == 8'hc7 | _GEN_2234; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2238 = i == 8'hc8 ? 1'h0 : i == 8'hc8 | _GEN_2236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2240 = i == 8'hc9 ? 1'h0 : i == 8'hc9 | _GEN_2238; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2241 = i == 8'h1 ? 1'h0 : _GEN_1913; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2242 = i == 8'h2 ? 1'h0 : _GEN_2241; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2243 = i == 8'h4 ? 1'h0 : _GEN_2242; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2244 = i == 8'h5 ? 1'h0 : _GEN_2243; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2245 = i == 8'ha ? 1'h0 : _GEN_2244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2246 = i == 8'h16 ? 1'h0 : _GEN_2245; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2247 = i == 8'h18 ? 1'h0 : _GEN_2246; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2248 = i == 8'h2e ? 1'h0 : _GEN_2247; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2249 = i == 8'h64 ? 1'h0 : _GEN_2248; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2250 = i == 8'hbd ? 1'h0 : _GEN_2249; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2251 = _GEN_3306 == 9'h17c ? 1'h0 : _GEN_2250; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2253 = _GEN_3306 == 9'h17d ? 1'h0 : _GEN_3306 == 9'h17c | _GEN_2251; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2255 = _GEN_3306 == 9'h17e ? 1'h0 : _GEN_3306 == 9'h17d | _GEN_2253; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2257 = _GEN_3306 == 9'h17f ? 1'h0 : _GEN_3306 == 9'h17e | _GEN_2255; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2259 = _GEN_3306 == 9'h180 ? 1'h0 : _GEN_3306 == 9'h17f | _GEN_2257; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2261 = _GEN_3306 == 9'h181 ? 1'h0 : _GEN_3306 == 9'h180 | _GEN_2259; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2263 = _GEN_3306 == 9'h182 ? 1'h0 : _GEN_3306 == 9'h181 | _GEN_2261; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2265 = _GEN_3306 == 9'h183 ? 1'h0 : _GEN_3306 == 9'h182 | _GEN_2263; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2267 = _GEN_3306 == 9'h184 ? 1'h0 : _GEN_3306 == 9'h183 | _GEN_2265; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2269 = _GEN_3306 == 9'h185 ? 1'h0 : _GEN_3306 == 9'h184 | _GEN_2267; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2271 = _GEN_3306 == 9'h186 ? 1'h0 : _GEN_3306 == 9'h185 | _GEN_2269; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2273 = _GEN_3306 == 9'h187 ? 1'h0 : _GEN_3306 == 9'h186 | _GEN_2271; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2275 = _GEN_3306 == 9'h188 ? 1'h0 : _GEN_3306 == 9'h187 | _GEN_2273; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2277 = _GEN_3306 == 9'h189 ? 1'h0 : _GEN_3306 == 9'h188 | _GEN_2275; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2279 = _GEN_3306 == 9'h18a ? 1'h0 : _GEN_3306 == 9'h189 | _GEN_2277; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2281 = _GEN_3306 == 9'h18b ? 1'h0 : _GEN_3306 == 9'h18a | _GEN_2279; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2283 = _GEN_3306 == 9'h18c ? 1'h0 : _GEN_3306 == 9'h18b | _GEN_2281; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2285 = _GEN_3306 == 9'h18d ? 1'h0 : _GEN_3306 == 9'h18c | _GEN_2283; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2287 = _GEN_3306 == 9'h18e ? 1'h0 : _GEN_3306 == 9'h18d | _GEN_2285; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2289 = _GEN_3306 == 9'h18f ? 1'h0 : _GEN_3306 == 9'h18e | _GEN_2287; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2291 = _GEN_3306 == 9'h190 ? 1'h0 : _GEN_3306 == 9'h18f | _GEN_2289; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2293 = _GEN_3306 == 9'h191 ? 1'h0 : _GEN_3306 == 9'h190 | _GEN_2291; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2295 = _GEN_3306 == 9'h192 ? 1'h0 : _GEN_3306 == 9'h191 | _GEN_2293; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2297 = _GEN_3306 == 9'h193 ? 1'h0 : _GEN_3306 == 9'h192 | _GEN_2295; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2299 = _GEN_3306 == 9'h194 ? 1'h0 : _GEN_3306 == 9'h193 | _GEN_2297; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2301 = i == 8'h1 ? 1'h0 : _GEN_3307 == 10'h311 | _GEN_2124; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2302 = i == 8'h2 ? 1'h0 : _GEN_2301; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2303 = i == 8'h4 ? 1'h0 : _GEN_2302; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2304 = i == 8'h5 ? 1'h0 : _GEN_2303; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2305 = i == 8'ha ? 1'h0 : _GEN_2304; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2306 = i == 8'h16 ? 1'h0 : _GEN_2305; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2307 = i == 8'h18 ? 1'h0 : _GEN_2306; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2308 = i == 8'h2e ? 1'h0 : _GEN_2307; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2309 = i == 8'h64 ? 1'h0 : _GEN_2308; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2310 = i == 8'hbd ? 1'h0 : _GEN_2309; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2311 = _GEN_3307 == 10'h2f9 ? 1'h0 : _GEN_2310; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2313 = _GEN_3307 == 10'h2fa ? 1'h0 : _GEN_3307 == 10'h2f9 | _GEN_2311; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2315 = _GEN_3307 == 10'h2fb ? 1'h0 : _GEN_3307 == 10'h2fa | _GEN_2313; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2317 = _GEN_3307 == 10'h2fc ? 1'h0 : _GEN_3307 == 10'h2fb | _GEN_2315; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2319 = _GEN_3307 == 10'h2fd ? 1'h0 : _GEN_3307 == 10'h2fc | _GEN_2317; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2321 = _GEN_3307 == 10'h2fe ? 1'h0 : _GEN_3307 == 10'h2fd | _GEN_2319; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2323 = _GEN_3307 == 10'h2ff ? 1'h0 : _GEN_3307 == 10'h2fe | _GEN_2321; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2325 = _GEN_3307 == 10'h300 ? 1'h0 : _GEN_3307 == 10'h2ff | _GEN_2323; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2327 = _GEN_3307 == 10'h301 ? 1'h0 : _GEN_3307 == 10'h300 | _GEN_2325; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2329 = _GEN_3307 == 10'h302 ? 1'h0 : _GEN_3307 == 10'h301 | _GEN_2327; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2331 = _GEN_3307 == 10'h303 ? 1'h0 : _GEN_3307 == 10'h302 | _GEN_2329; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2333 = _GEN_3307 == 10'h304 ? 1'h0 : _GEN_3307 == 10'h303 | _GEN_2331; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2335 = _GEN_3307 == 10'h305 ? 1'h0 : _GEN_3307 == 10'h304 | _GEN_2333; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2337 = _GEN_3307 == 10'h306 ? 1'h0 : _GEN_3307 == 10'h305 | _GEN_2335; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2339 = _GEN_3307 == 10'h307 ? 1'h0 : _GEN_3307 == 10'h306 | _GEN_2337; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2341 = _GEN_3307 == 10'h308 ? 1'h0 : _GEN_3307 == 10'h307 | _GEN_2339; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2343 = _GEN_3307 == 10'h309 ? 1'h0 : _GEN_3307 == 10'h308 | _GEN_2341; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2345 = _GEN_3307 == 10'h30a ? 1'h0 : _GEN_3307 == 10'h309 | _GEN_2343; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2347 = _GEN_3307 == 10'h30b ? 1'h0 : _GEN_3307 == 10'h30a | _GEN_2345; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2349 = _GEN_3307 == 10'h30c ? 1'h0 : _GEN_3307 == 10'h30b | _GEN_2347; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2351 = _GEN_3307 == 10'h30d ? 1'h0 : _GEN_3307 == 10'h30c | _GEN_2349; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2353 = _GEN_3307 == 10'h30e ? 1'h0 : _GEN_3307 == 10'h30d | _GEN_2351; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2355 = _GEN_3307 == 10'h30f ? 1'h0 : _GEN_3307 == 10'h30e | _GEN_2353; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2357 = _GEN_3307 == 10'h310 ? 1'h0 : _GEN_3307 == 10'h30f | _GEN_2355; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2359 = _GEN_3307 == 10'h311 ? 1'h0 : _GEN_3307 == 10'h310 | _GEN_2357; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2361 = _GEN_3307 == 10'h312 ? 1'h0 : _GEN_3307 == 10'h311 | _GEN_2359; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2363 = _GEN_3307 == 10'h313 ? 1'h0 : _GEN_3307 == 10'h312 | _GEN_2361; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2365 = _GEN_3307 == 10'h314 ? 1'h0 : _GEN_3307 == 10'h313 | _GEN_2363; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2367 = _GEN_3307 == 10'h315 ? 1'h0 : _GEN_3307 == 10'h314 | _GEN_2365; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2369 = _GEN_3307 == 10'h316 ? 1'h0 : _GEN_3307 == 10'h315 | _GEN_2367; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2371 = _GEN_3307 == 10'h317 ? 1'h0 : _GEN_3307 == 10'h316 | _GEN_2369; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2373 = _GEN_3307 == 10'h318 ? 1'h0 : _GEN_3307 == 10'h317 | _GEN_2371; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2375 = _GEN_3307 == 10'h319 ? 1'h0 : _GEN_3307 == 10'h318 | _GEN_2373; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2377 = _GEN_3307 == 10'h31a ? 1'h0 : _GEN_3307 == 10'h319 | _GEN_2375; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2379 = _GEN_3307 == 10'h31b ? 1'h0 : _GEN_3307 == 10'h31a | _GEN_2377; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2381 = _GEN_3307 == 10'h31c ? 1'h0 : _GEN_3307 == 10'h31b | _GEN_2379; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2383 = _GEN_3307 == 10'h31d ? 1'h0 : _GEN_3307 == 10'h31c | _GEN_2381; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2385 = _GEN_3307 == 10'h31e ? 1'h0 : _GEN_3307 == 10'h31d | _GEN_2383; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2387 = _GEN_3307 == 10'h31f ? 1'h0 : _GEN_3307 == 10'h31e | _GEN_2385; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2389 = _GEN_3307 == 10'h320 ? 1'h0 : _GEN_3307 == 10'h31f | _GEN_2387; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2391 = _GEN_3307 == 10'h321 ? 1'h0 : _GEN_3307 == 10'h320 | _GEN_2389; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2393 = _GEN_3307 == 10'h322 ? 1'h0 : _GEN_3307 == 10'h321 | _GEN_2391; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2395 = _GEN_3307 == 10'h323 ? 1'h0 : _GEN_3307 == 10'h322 | _GEN_2393; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2397 = _GEN_3307 == 10'h324 ? 1'h0 : _GEN_3307 == 10'h323 | _GEN_2395; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2399 = _GEN_3307 == 10'h325 ? 1'h0 : _GEN_3307 == 10'h324 | _GEN_2397; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2401 = _GEN_3307 == 10'h326 ? 1'h0 : _GEN_3307 == 10'h325 | _GEN_2399; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2403 = _GEN_3307 == 10'h327 ? 1'h0 : _GEN_3307 == 10'h326 | _GEN_2401; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2405 = _GEN_3307 == 10'h328 ? 1'h0 : _GEN_3307 == 10'h327 | _GEN_2403; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2407 = _GEN_3307 == 10'h329 ? 1'h0 : _GEN_3307 == 10'h328 | _GEN_2405; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2409 = _GEN_3307 == 10'h32a ? 1'h0 : _GEN_3307 == 10'h329 | _GEN_2407; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2411 = i == 8'h0 ? 1'h0 : i == 8'hc5 | _GEN_2133; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2412 = i == 8'h1 ? 1'h0 : _GEN_2411; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2413 = i == 8'h3 ? 1'h0 : _GEN_2412; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2417 = i == 8'h22 ? 1'h0 : i == 8'h22 | (i == 8'h10 | (i == 8'h7 | _GEN_2413)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2418 = i == 8'h0 ? 1'h0 : i == 8'hc9 | _GEN_2149; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2419 = i == 8'h1 ? 1'h0 : _GEN_2418; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2421 = i == 8'h8 ? 1'h0 : i == 8'h7 | _GEN_2419; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2422 = i == 8'h11 ? 1'h0 : _GEN_2421; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2424 = i == 8'h22 ? 1'h0 : i == 8'h21 | _GEN_2422; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2426 = i == 8'h23 ? 1'h0 : i == 8'h22 | _GEN_2424; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2427 = i == 8'h44 ? 1'h0 : _GEN_2426; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2429 = i == 8'h47 ? 1'h0 : i == 8'h47 | _GEN_2427; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2431 = i == 8'h89 ? 1'h0 : i == 8'h89 | _GEN_2429; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2432 = i == 8'h0 ? 1'h0 : _GEN_2172; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2433 = i == 8'h1 ? 1'h0 : _GEN_2432; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2434 = i == 8'h7 ? 1'h0 : _GEN_2433; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2435 = i == 8'h8 ? 1'h0 : _GEN_2434; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2436 = i == 8'h11 ? 1'h0 : _GEN_2435; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2437 = i == 8'h21 ? 1'h0 : _GEN_2436; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2439 = i == 8'h45 ? 1'h0 : i == 8'h44 | _GEN_2437; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2441 = i == 8'h47 ? 1'h0 : i == 8'h46 | _GEN_2439; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2443 = i == 8'h48 ? 1'h0 : i == 8'h47 | _GEN_2441; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2444 = i == 8'h89 ? 1'h0 : _GEN_2443; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2447 = i == 8'h8b ? 1'h0 : i == 8'h8b | (i == 8'h89 | _GEN_2444); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2449 = i == 8'h8e ? 1'h0 : i == 8'h8e | _GEN_2447; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2451 = i == 8'h91 ? 1'h0 : i == 8'h91 | _GEN_2449; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2452 = i == 8'h0 ? 1'h0 : _GEN_2206; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2453 = i == 8'h1 ? 1'h0 : _GEN_2452; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2454 = i == 8'h7 ? 1'h0 : _GEN_2453; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2455 = i == 8'h8 ? 1'h0 : _GEN_2454; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2456 = i == 8'h11 ? 1'h0 : _GEN_2455; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2457 = i == 8'h21 ? 1'h0 : _GEN_2456; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2458 = i == 8'h45 ? 1'h0 : _GEN_2457; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2460 = i == 8'h89 ? 1'h0 : i == 8'h47 | _GEN_2458; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2463 = i == 8'h8a ? 1'h0 : i == 8'h8a | (i == 8'h89 | _GEN_2460); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2464 = i == 8'h8b ? 1'h0 : _GEN_2463; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2467 = i == 8'h8d ? 1'h0 : i == 8'h8d | (i == 8'h8b | _GEN_2464); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2468 = i == 8'h8e ? 1'h0 : _GEN_2467; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2471 = i == 8'h8f ? 1'h0 : i == 8'h8f | (i == 8'h8e | _GEN_2468); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2472 = i == 8'h91 ? 1'h0 : _GEN_2471; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2475 = i == 8'h92 ? 1'h0 : i == 8'h92 | (i == 8'h91 | _GEN_2472); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2476 = i == 8'h0 ? 1'h0 : _GEN_2240; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2477 = i == 8'h1 ? 1'h0 : _GEN_2476; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2479 = i == 8'h8 ? 1'h0 : i == 8'h7 | _GEN_2477; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2480 = i == 8'h11 ? 1'h0 : _GEN_2479; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2483 = i == 8'h45 ? 1'h0 : i == 8'h44 | (i == 8'h21 | _GEN_2480); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2485 = i == 8'h47 ? 1'h0 : i == 8'h46 | _GEN_2483; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2487 = i == 8'h8a ? 1'h0 : i == 8'h48 | _GEN_2485; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2490 = i == 8'h8c ? 1'h0 : i == 8'h8c | (i == 8'h8a | _GEN_2487); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2491 = i == 8'h8e ? 1'h0 : _GEN_2490; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2494 = i == 8'h90 ? 1'h0 : i == 8'h90 | (i == 8'h8e | _GEN_2491); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2495 = i == 8'h92 ? 1'h0 : _GEN_2494; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2497 = i == 8'h0 ? 1'h0 : _GEN_3306 == 9'h194 | _GEN_2299; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2498 = i == 8'h1 ? 1'h0 : _GEN_2497; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2499 = i == 8'h7 ? 1'h0 : _GEN_2498; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2500 = i == 8'h8 ? 1'h0 : _GEN_2499; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2501 = i == 8'h11 ? 1'h0 : _GEN_2500; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2502 = i == 8'h21 ? 1'h0 : _GEN_2501; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2503 = i == 8'h89 ? 1'h0 : _GEN_2502; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2506 = i == 8'h8a ? 1'h0 : i == 8'h8a | (i == 8'h89 | _GEN_2503); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2507 = i == 8'h8b ? 1'h0 : _GEN_2506; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2510 = i == 8'h8c ? 1'h0 : i == 8'h8c | (i == 8'h8b | _GEN_2507); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2511 = i == 8'h8d ? 1'h0 : _GEN_2510; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2514 = i == 8'h8e ? 1'h0 : i == 8'h8e | (i == 8'h8d | _GEN_2511); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2515 = i == 8'h8f ? 1'h0 : _GEN_2514; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2518 = i == 8'h90 ? 1'h0 : i == 8'h90 | (i == 8'h8f | _GEN_2515); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2519 = i == 8'h91 ? 1'h0 : _GEN_2518; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2522 = i == 8'h92 ? 1'h0 : i == 8'h92 | (i == 8'h91 | _GEN_2519); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2523 = i == 8'h0 ? 1'h0 : _GEN_3307 == 10'h32a | _GEN_2409; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2524 = i == 8'h1 ? 1'h0 : _GEN_2523; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2525 = i == 8'h7 ? 1'h0 : _GEN_2524; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2526 = i == 8'h8 ? 1'h0 : _GEN_2525; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2527 = i == 8'h11 ? 1'h0 : _GEN_2526; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2528 = i == 8'h21 ? 1'h0 : _GEN_2527; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2529 = i == 8'h89 ? 1'h0 : _GEN_2528; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2531 = i == 8'h8a ? 1'h0 : i == 8'h89 | _GEN_2529; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2533 = i == 8'h8b ? 1'h0 : i == 8'h8a | _GEN_2531; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2535 = i == 8'h8c ? 1'h0 : i == 8'h8b | _GEN_2533; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2537 = i == 8'h8d ? 1'h0 : i == 8'h8c | _GEN_2535; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2539 = i == 8'h8e ? 1'h0 : i == 8'h8d | _GEN_2537; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2541 = i == 8'h8f ? 1'h0 : i == 8'h8e | _GEN_2539; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2543 = i == 8'h90 ? 1'h0 : i == 8'h8f | _GEN_2541; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2545 = i == 8'h91 ? 1'h0 : i == 8'h90 | _GEN_2543; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2547 = i == 8'h92 ? 1'h0 : i == 8'h91 | _GEN_2545; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2549 = i == 8'h0 ? 1'h0 : _GEN_2417; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2550 = i == 8'h3 ? 1'h0 : _GEN_2549; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2551 = i == 8'h4 ? 1'h0 : _GEN_2550; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2553 = i == 8'h9 ? 1'h0 : i == 8'h8 | _GEN_2551; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2555 = i == 8'h13 ? 1'h0 : i == 8'h11 | _GEN_2553; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2558 = i == 8'h27 ? 1'h0 : i == 8'h27 | (i == 8'h23 | _GEN_2555); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2560 = i == 8'h8f ? 1'h0 : i == 8'h47 | _GEN_2558; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2562 = i == 8'h0 ? 1'h0 : _GEN_2431; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2563 = i == 8'h4 ? 1'h0 : _GEN_2562; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2564 = i == 8'h7 ? 1'h0 : _GEN_2563; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2565 = i == 8'h9 ? 1'h0 : _GEN_2564; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2566 = i == 8'h10 ? 1'h0 : _GEN_2565; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2570 = i == 8'h23 ? 1'h0 : i == 8'h22 | (i == 8'h12 | (i == 8'h11 | _GEN_2566)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2572 = i == 8'h27 ? 1'h0 : i == 8'h26 | _GEN_2570; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2574 = i == 8'h28 ? 1'h0 : i == 8'h27 | _GEN_2572; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2575 = i == 8'h45 ? 1'h0 : _GEN_2574; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2576 = i == 8'h47 ? 1'h0 : _GEN_2575; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2577 = i == 8'h4e ? 1'h0 : _GEN_2576; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2579 = i == 8'h51 ? 1'h0 : i == 8'h51 | _GEN_2577; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2580 = i == 8'h8c ? 1'h0 : _GEN_2579; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2583 = i == 8'h8f ? 1'h0 : i == 8'h8f | (i == 8'h8c | _GEN_2580); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2585 = i == 8'h9d ? 1'h0 : i == 8'h9d | _GEN_2583; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2586 = i == 8'h0 ? 1'h0 : _GEN_2451; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2587 = i == 8'h4 ? 1'h0 : _GEN_2586; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2588 = i == 8'h7 ? 1'h0 : _GEN_2587; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2589 = i == 8'h9 ? 1'h0 : _GEN_2588; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2590 = i == 8'h10 ? 1'h0 : _GEN_2589; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2591 = i == 8'h11 ? 1'h0 : _GEN_2590; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2592 = i == 8'h12 ? 1'h0 : _GEN_2591; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2594 = i == 8'h26 ? 1'h0 : i == 8'h23 | _GEN_2592; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2596 = i == 8'h46 ? 1'h0 : i == 8'h45 | _GEN_2594; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2598 = i == 8'h47 ? 1'h0 : i == 8'h46 | _GEN_2596; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2600 = i == 8'h4f ? 1'h0 : i == 8'h4e | _GEN_2598; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2602 = i == 8'h51 ? 1'h0 : i == 8'h50 | _GEN_2600; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2604 = i == 8'h52 ? 1'h0 : i == 8'h51 | _GEN_2602; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2606 = i == 8'h8c ? 1'h0 : i == 8'h8c | _GEN_2604; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2608 = i == 8'h8f ? 1'h0 : i == 8'h8f | _GEN_2606; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2609 = i == 8'h9d ? 1'h0 : _GEN_2608; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2612 = i == 8'h9f ? 1'h0 : i == 8'h9f | (i == 8'h9d | _GEN_2609); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2614 = i == 8'ha2 ? 1'h0 : i == 8'ha2 | _GEN_2612; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2616 = i == 8'ha5 ? 1'h0 : i == 8'ha5 | _GEN_2614; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2617 = i == 8'h0 ? 1'h0 : _GEN_2475; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2618 = i == 8'h4 ? 1'h0 : _GEN_2617; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2619 = i == 8'h7 ? 1'h0 : _GEN_2618; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2620 = i == 8'h9 ? 1'h0 : _GEN_2619; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2621 = i == 8'h11 ? 1'h0 : _GEN_2620; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2622 = i == 8'h12 ? 1'h0 : _GEN_2621; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2623 = i == 8'h21 ? 1'h0 : _GEN_2622; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2624 = i == 8'h26 ? 1'h0 : _GEN_2623; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2625 = i == 8'h44 ? 1'h0 : _GEN_2624; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2628 = i == 8'h46 ? 1'h0 : i == 8'h46 | (i == 8'h44 | _GEN_2625); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2629 = i == 8'h48 ? 1'h0 : _GEN_2628; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2631 = i == 8'h4f ? 1'h0 : i == 8'h48 | _GEN_2629; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2633 = i == 8'h8b ? 1'h0 : i == 8'h51 | _GEN_2631; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2636 = i == 8'h8c ? 1'h0 : i == 8'h8c | (i == 8'h8b | _GEN_2633); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2638 = i == 8'h8f ? 1'h0 : i == 8'h8f | _GEN_2636; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2639 = i == 8'h90 ? 1'h0 : _GEN_2638; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2641 = i == 8'h9d ? 1'h0 : i == 8'h90 | _GEN_2639; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2644 = i == 8'h9e ? 1'h0 : i == 8'h9e | (i == 8'h9d | _GEN_2641); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2645 = i == 8'h9f ? 1'h0 : _GEN_2644; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2648 = i == 8'ha1 ? 1'h0 : i == 8'ha1 | (i == 8'h9f | _GEN_2645); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2649 = i == 8'ha2 ? 1'h0 : _GEN_2648; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2652 = i == 8'ha3 ? 1'h0 : i == 8'ha3 | (i == 8'ha2 | _GEN_2649); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2653 = i == 8'ha5 ? 1'h0 : _GEN_2652; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2656 = i == 8'ha6 ? 1'h0 : i == 8'ha6 | (i == 8'ha5 | _GEN_2653); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2657 = i == 8'h0 ? 1'h0 : i == 8'h92 | _GEN_2495; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2658 = i == 8'h4 ? 1'h0 : _GEN_2657; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2659 = i == 8'h7 ? 1'h0 : _GEN_2658; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2660 = i == 8'h9 ? 1'h0 : _GEN_2659; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2663 = i == 8'h21 ? 1'h0 : i == 8'h12 | (i == 8'h11 | _GEN_2660); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2666 = i == 8'h4f ? 1'h0 : i == 8'h4e | (i == 8'h26 | _GEN_2663); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2668 = i == 8'h51 ? 1'h0 : i == 8'h50 | _GEN_2666; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2670 = i == 8'h89 ? 1'h0 : i == 8'h52 | _GEN_2668; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2672 = i == 8'h8a ? 1'h0 : i == 8'h89 | _GEN_2670; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2675 = i == 8'h8b ? 1'h0 : i == 8'h8b | (i == 8'h8a | _GEN_2672); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2677 = i == 8'h8c ? 1'h0 : i == 8'h8c | _GEN_2675; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2678 = i == 8'h8d ? 1'h0 : _GEN_2677; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2680 = i == 8'h8e ? 1'h0 : i == 8'h8d | _GEN_2678; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2683 = i == 8'h8f ? 1'h0 : i == 8'h8f | (i == 8'h8e | _GEN_2680); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2685 = i == 8'h90 ? 1'h0 : i == 8'h90 | _GEN_2683; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2686 = i == 8'h91 ? 1'h0 : _GEN_2685; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2688 = i == 8'h92 ? 1'h0 : i == 8'h91 | _GEN_2686; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2690 = i == 8'h9e ? 1'h0 : i == 8'h92 | _GEN_2688; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2693 = i == 8'ha0 ? 1'h0 : i == 8'ha0 | (i == 8'h9e | _GEN_2690); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2694 = i == 8'ha2 ? 1'h0 : _GEN_2693; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2697 = i == 8'ha4 ? 1'h0 : i == 8'ha4 | (i == 8'ha2 | _GEN_2694); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2698 = i == 8'ha6 ? 1'h0 : _GEN_2697; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2700 = i == 8'h0 ? 1'h0 : _GEN_2522; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2701 = i == 8'h4 ? 1'h0 : _GEN_2700; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2702 = i == 8'h7 ? 1'h0 : _GEN_2701; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2703 = i == 8'h9 ? 1'h0 : _GEN_2702; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2704 = i == 8'h11 ? 1'h0 : _GEN_2703; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2705 = i == 8'h12 ? 1'h0 : _GEN_2704; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2706 = i == 8'h21 ? 1'h0 : _GEN_2705; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2707 = i == 8'h26 ? 1'h0 : _GEN_2706; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2708 = i == 8'h44 ? 1'h0 : _GEN_2707; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2710 = i == 8'h45 ? 1'h0 : i == 8'h44 | _GEN_2708; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2712 = i == 8'h46 ? 1'h0 : i == 8'h45 | _GEN_2710; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2714 = i == 8'h47 ? 1'h0 : i == 8'h46 | _GEN_2712; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2716 = i == 8'h48 ? 1'h0 : i == 8'h47 | _GEN_2714; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2718 = i == 8'h9d ? 1'h0 : i == 8'h48 | _GEN_2716; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2721 = i == 8'h9e ? 1'h0 : i == 8'h9e | (i == 8'h9d | _GEN_2718); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2722 = i == 8'h9f ? 1'h0 : _GEN_2721; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2725 = i == 8'ha0 ? 1'h0 : i == 8'ha0 | (i == 8'h9f | _GEN_2722); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2726 = i == 8'ha1 ? 1'h0 : _GEN_2725; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2729 = i == 8'ha2 ? 1'h0 : i == 8'ha2 | (i == 8'ha1 | _GEN_2726); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2730 = i == 8'ha3 ? 1'h0 : _GEN_2729; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2733 = i == 8'ha4 ? 1'h0 : i == 8'ha4 | (i == 8'ha3 | _GEN_2730); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2734 = i == 8'ha5 ? 1'h0 : _GEN_2733; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2737 = i == 8'ha6 ? 1'h0 : i == 8'ha6 | (i == 8'ha5 | _GEN_2734); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2738 = i == 8'h0 ? 1'h0 : i == 8'h92 | _GEN_2547; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2739 = i == 8'h4 ? 1'h0 : _GEN_2738; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2740 = i == 8'h7 ? 1'h0 : _GEN_2739; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2741 = i == 8'h9 ? 1'h0 : _GEN_2740; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2742 = i == 8'h11 ? 1'h0 : _GEN_2741; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2743 = i == 8'h12 ? 1'h0 : _GEN_2742; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2744 = i == 8'h21 ? 1'h0 : _GEN_2743; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2745 = i == 8'h26 ? 1'h0 : _GEN_2744; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2746 = i == 8'h89 ? 1'h0 : _GEN_2745; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2748 = i == 8'h8a ? 1'h0 : i == 8'h89 | _GEN_2746; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2750 = i == 8'h8b ? 1'h0 : i == 8'h8a | _GEN_2748; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2752 = i == 8'h8c ? 1'h0 : i == 8'h8b | _GEN_2750; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2754 = i == 8'h8d ? 1'h0 : i == 8'h8c | _GEN_2752; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2756 = i == 8'h8e ? 1'h0 : i == 8'h8d | _GEN_2754; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2758 = i == 8'h8f ? 1'h0 : i == 8'h8e | _GEN_2756; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2760 = i == 8'h90 ? 1'h0 : i == 8'h8f | _GEN_2758; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2762 = i == 8'h91 ? 1'h0 : i == 8'h90 | _GEN_2760; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2764 = i == 8'h92 ? 1'h0 : i == 8'h91 | _GEN_2762; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2766 = i == 8'h9d ? 1'h0 : i == 8'h92 | _GEN_2764; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2768 = i == 8'h9e ? 1'h0 : i == 8'h9d | _GEN_2766; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2770 = i == 8'h9f ? 1'h0 : i == 8'h9e | _GEN_2768; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2772 = i == 8'ha0 ? 1'h0 : i == 8'h9f | _GEN_2770; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2774 = i == 8'ha1 ? 1'h0 : i == 8'ha0 | _GEN_2772; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2776 = i == 8'ha2 ? 1'h0 : i == 8'ha1 | _GEN_2774; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2778 = i == 8'ha3 ? 1'h0 : i == 8'ha2 | _GEN_2776; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2780 = i == 8'ha4 ? 1'h0 : i == 8'ha3 | _GEN_2778; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2782 = i == 8'ha5 ? 1'h0 : i == 8'ha4 | _GEN_2780; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2784 = i == 8'ha6 ? 1'h0 : i == 8'ha5 | _GEN_2782; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2786 = i == 8'h0 ? 1'h0 : i == 8'h8f | _GEN_2560; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2787 = i == 8'h1 ? 1'h0 : _GEN_2786; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2789 = i == 8'ha ? 1'h0 : i == 8'h9 | _GEN_2787; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2790 = i == 8'h13 ? 1'h0 : _GEN_2789; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2794 = i == 8'h2c ? 1'h0 : i == 8'h2c | (i == 8'h28 | (i == 8'h15 | _GEN_2790)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2796 = i == 8'ha3 ? 1'h0 : i == 8'h51 | _GEN_2794; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2798 = i == 8'h0 ? 1'h0 : _GEN_2585; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2799 = i == 8'h1 ? 1'h0 : _GEN_2798; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2801 = i == 8'h16 ? 1'h0 : i == 8'h9 | _GEN_2799; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2803 = i == 8'h28 ? 1'h0 : i == 8'h27 | _GEN_2801; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2805 = i == 8'h2c ? 1'h0 : i == 8'h2b | _GEN_2803; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2807 = i == 8'h2d ? 1'h0 : i == 8'h2c | _GEN_2805; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2808 = i == 8'h4f ? 1'h0 : _GEN_2807; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2809 = i == 8'h51 ? 1'h0 : _GEN_2808; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2810 = i == 8'h58 ? 1'h0 : _GEN_2809; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2812 = i == 8'h5b ? 1'h0 : i == 8'h5b | _GEN_2810; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2813 = i == 8'ha0 ? 1'h0 : _GEN_2812; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2816 = i == 8'ha3 ? 1'h0 : i == 8'ha3 | (i == 8'ha0 | _GEN_2813); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2818 = i == 8'hb1 ? 1'h0 : i == 8'hb1 | _GEN_2816; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2819 = i == 8'h0 ? 1'h0 : _GEN_2616; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2820 = i == 8'h1 ? 1'h0 : _GEN_2819; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2821 = i == 8'h9 ? 1'h0 : _GEN_2820; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2822 = i == 8'h16 ? 1'h0 : _GEN_2821; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2824 = i == 8'h2b ? 1'h0 : i == 8'h28 | _GEN_2822; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2826 = i == 8'h50 ? 1'h0 : i == 8'h4f | _GEN_2824; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2828 = i == 8'h51 ? 1'h0 : i == 8'h50 | _GEN_2826; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2830 = i == 8'h59 ? 1'h0 : i == 8'h58 | _GEN_2828; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2832 = i == 8'h5b ? 1'h0 : i == 8'h5a | _GEN_2830; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2834 = i == 8'h5c ? 1'h0 : i == 8'h5b | _GEN_2832; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2836 = i == 8'ha0 ? 1'h0 : i == 8'ha0 | _GEN_2834; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2838 = i == 8'ha3 ? 1'h0 : i == 8'ha3 | _GEN_2836; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2839 = i == 8'hb1 ? 1'h0 : _GEN_2838; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2842 = i == 8'hb3 ? 1'h0 : i == 8'hb3 | (i == 8'hb1 | _GEN_2839); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2844 = i == 8'hb6 ? 1'h0 : i == 8'hb6 | _GEN_2842; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2846 = i == 8'hb9 ? 1'h0 : i == 8'hb9 | _GEN_2844; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2847 = i == 8'h0 ? 1'h0 : _GEN_2656; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2848 = i == 8'h3 ? 1'h0 : _GEN_2847; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2849 = i == 8'h8 ? 1'h0 : _GEN_2848; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2850 = i == 8'h9 ? 1'h0 : _GEN_2849; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2851 = i == 8'h12 ? 1'h0 : _GEN_2850; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2852 = i == 8'h16 ? 1'h0 : _GEN_2851; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2853 = i == 8'h26 ? 1'h0 : _GEN_2852; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2854 = i == 8'h2b ? 1'h0 : _GEN_2853; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2855 = i == 8'h4e ? 1'h0 : _GEN_2854; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2858 = i == 8'h50 ? 1'h0 : i == 8'h50 | (i == 8'h4e | _GEN_2855); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2859 = i == 8'h52 ? 1'h0 : _GEN_2858; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2861 = i == 8'h59 ? 1'h0 : i == 8'h52 | _GEN_2859; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2863 = i == 8'h9f ? 1'h0 : i == 8'h5b | _GEN_2861; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2866 = i == 8'ha0 ? 1'h0 : i == 8'ha0 | (i == 8'h9f | _GEN_2863); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2868 = i == 8'ha3 ? 1'h0 : i == 8'ha3 | _GEN_2866; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2869 = i == 8'ha4 ? 1'h0 : _GEN_2868; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2871 = i == 8'hb1 ? 1'h0 : i == 8'ha4 | _GEN_2869; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2874 = i == 8'hb2 ? 1'h0 : i == 8'hb2 | (i == 8'hb1 | _GEN_2871); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2875 = i == 8'hb3 ? 1'h0 : _GEN_2874; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2878 = i == 8'hb5 ? 1'h0 : i == 8'hb5 | (i == 8'hb3 | _GEN_2875); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2879 = i == 8'hb6 ? 1'h0 : _GEN_2878; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2882 = i == 8'hb7 ? 1'h0 : i == 8'hb7 | (i == 8'hb6 | _GEN_2879); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2883 = i == 8'hb9 ? 1'h0 : _GEN_2882; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2886 = i == 8'hba ? 1'h0 : i == 8'hba | (i == 8'hb9 | _GEN_2883); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2887 = i == 8'h0 ? 1'h0 : i == 8'ha6 | _GEN_2698; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2888 = i == 8'h3 ? 1'h0 : _GEN_2887; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2889 = i == 8'h8 ? 1'h0 : _GEN_2888; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2891 = i == 8'h12 ? 1'h0 : i == 8'h9 | _GEN_2889; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2892 = i == 8'h16 ? 1'h0 : _GEN_2891; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2893 = i == 8'h26 ? 1'h0 : _GEN_2892; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2896 = i == 8'h59 ? 1'h0 : i == 8'h58 | (i == 8'h2b | _GEN_2893); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2898 = i == 8'h5b ? 1'h0 : i == 8'h5a | _GEN_2896; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2900 = i == 8'h9d ? 1'h0 : i == 8'h5c | _GEN_2898; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2902 = i == 8'h9e ? 1'h0 : i == 8'h9d | _GEN_2900; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2905 = i == 8'h9f ? 1'h0 : i == 8'h9f | (i == 8'h9e | _GEN_2902); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2907 = i == 8'ha0 ? 1'h0 : i == 8'ha0 | _GEN_2905; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2908 = i == 8'ha1 ? 1'h0 : _GEN_2907; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2910 = i == 8'ha2 ? 1'h0 : i == 8'ha1 | _GEN_2908; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2913 = i == 8'ha3 ? 1'h0 : i == 8'ha3 | (i == 8'ha2 | _GEN_2910); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2915 = i == 8'ha4 ? 1'h0 : i == 8'ha4 | _GEN_2913; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2916 = i == 8'ha5 ? 1'h0 : _GEN_2915; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2918 = i == 8'ha6 ? 1'h0 : i == 8'ha5 | _GEN_2916; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2920 = i == 8'hb2 ? 1'h0 : i == 8'ha6 | _GEN_2918; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2923 = i == 8'hb4 ? 1'h0 : i == 8'hb4 | (i == 8'hb2 | _GEN_2920); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2924 = i == 8'hb6 ? 1'h0 : _GEN_2923; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2927 = i == 8'hb8 ? 1'h0 : i == 8'hb8 | (i == 8'hb6 | _GEN_2924); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2928 = i == 8'hba ? 1'h0 : _GEN_2927; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2930 = i == 8'h0 ? 1'h0 : _GEN_2737; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2931 = i == 8'h3 ? 1'h0 : _GEN_2930; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2932 = i == 8'h8 ? 1'h0 : _GEN_2931; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2933 = i == 8'h9 ? 1'h0 : _GEN_2932; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2934 = i == 8'h12 ? 1'h0 : _GEN_2933; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2935 = i == 8'h16 ? 1'h0 : _GEN_2934; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2936 = i == 8'h26 ? 1'h0 : _GEN_2935; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2937 = i == 8'h2b ? 1'h0 : _GEN_2936; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2938 = i == 8'h4e ? 1'h0 : _GEN_2937; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2940 = i == 8'h4f ? 1'h0 : i == 8'h4e | _GEN_2938; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2942 = i == 8'h50 ? 1'h0 : i == 8'h4f | _GEN_2940; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2944 = i == 8'h51 ? 1'h0 : i == 8'h50 | _GEN_2942; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2946 = i == 8'h52 ? 1'h0 : i == 8'h51 | _GEN_2944; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2948 = i == 8'hb1 ? 1'h0 : i == 8'h52 | _GEN_2946; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2951 = i == 8'hb2 ? 1'h0 : i == 8'hb2 | (i == 8'hb1 | _GEN_2948); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2952 = i == 8'hb3 ? 1'h0 : _GEN_2951; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2955 = i == 8'hb4 ? 1'h0 : i == 8'hb4 | (i == 8'hb3 | _GEN_2952); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2956 = i == 8'hb5 ? 1'h0 : _GEN_2955; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2959 = i == 8'hb6 ? 1'h0 : i == 8'hb6 | (i == 8'hb5 | _GEN_2956); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2960 = i == 8'hb7 ? 1'h0 : _GEN_2959; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2963 = i == 8'hb8 ? 1'h0 : i == 8'hb8 | (i == 8'hb7 | _GEN_2960); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2964 = i == 8'hb9 ? 1'h0 : _GEN_2963; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2967 = i == 8'hba ? 1'h0 : i == 8'hba | (i == 8'hb9 | _GEN_2964); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2968 = i == 8'h0 ? 1'h0 : i == 8'ha6 | _GEN_2784; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2969 = i == 8'h3 ? 1'h0 : _GEN_2968; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2970 = i == 8'h8 ? 1'h0 : _GEN_2969; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2971 = i == 8'h9 ? 1'h0 : _GEN_2970; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2972 = i == 8'h12 ? 1'h0 : _GEN_2971; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2973 = i == 8'h16 ? 1'h0 : _GEN_2972; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2974 = i == 8'h26 ? 1'h0 : _GEN_2973; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2975 = i == 8'h2b ? 1'h0 : _GEN_2974; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2976 = i == 8'h9d ? 1'h0 : _GEN_2975; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2978 = i == 8'h9e ? 1'h0 : i == 8'h9d | _GEN_2976; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2980 = i == 8'h9f ? 1'h0 : i == 8'h9e | _GEN_2978; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2982 = i == 8'ha0 ? 1'h0 : i == 8'h9f | _GEN_2980; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2984 = i == 8'ha1 ? 1'h0 : i == 8'ha0 | _GEN_2982; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2986 = i == 8'ha2 ? 1'h0 : i == 8'ha1 | _GEN_2984; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2988 = i == 8'ha3 ? 1'h0 : i == 8'ha2 | _GEN_2986; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2990 = i == 8'ha4 ? 1'h0 : i == 8'ha3 | _GEN_2988; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2992 = i == 8'ha5 ? 1'h0 : i == 8'ha4 | _GEN_2990; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2994 = i == 8'ha6 ? 1'h0 : i == 8'ha5 | _GEN_2992; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2996 = i == 8'hb1 ? 1'h0 : i == 8'ha6 | _GEN_2994; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_2998 = i == 8'hb2 ? 1'h0 : i == 8'hb1 | _GEN_2996; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3000 = i == 8'hb3 ? 1'h0 : i == 8'hb2 | _GEN_2998; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3002 = i == 8'hb4 ? 1'h0 : i == 8'hb3 | _GEN_3000; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3004 = i == 8'hb5 ? 1'h0 : i == 8'hb4 | _GEN_3002; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3006 = i == 8'hb6 ? 1'h0 : i == 8'hb5 | _GEN_3004; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3008 = i == 8'hb7 ? 1'h0 : i == 8'hb6 | _GEN_3006; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3010 = i == 8'hb8 ? 1'h0 : i == 8'hb7 | _GEN_3008; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3012 = i == 8'hb9 ? 1'h0 : i == 8'hb8 | _GEN_3010; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3014 = i == 8'hba ? 1'h0 : i == 8'hb9 | _GEN_3012; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3016 = i == 8'h1 ? 1'h0 : i == 8'ha3 | _GEN_2796; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3017 = i == 8'h2 ? 1'h0 : _GEN_3016; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3018 = i == 8'h4 ? 1'h0 : _GEN_3017; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3019 = i == 8'h5 ? 1'h0 : _GEN_3018; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3020 = i == 8'ha ? 1'h0 : _GEN_3019; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3023 = i == 8'h18 ? 1'h0 : i == 8'h16 | (i == 8'hb | _GEN_3020); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3026 = i == 8'h31 ? 1'h0 : i == 8'h31 | (i == 8'h2d | _GEN_3023); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3028 = i == 8'hb7 ? 1'h0 : i == 8'h5b | _GEN_3026; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3029 = i == 8'hb7 | _GEN_3028; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3030 = i == 8'h1 ? 1'h0 : _GEN_2818; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3031 = i == 8'h2 ? 1'h0 : _GEN_3030; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3032 = i == 8'h4 ? 1'h0 : _GEN_3031; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3033 = i == 8'h5 ? 1'h0 : _GEN_3032; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3034 = i == 8'h15 ? 1'h0 : _GEN_3033; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3038 = i == 8'h2d ? 1'h0 : i == 8'h2c | (i == 8'h17 | (i == 8'h16 | _GEN_3034)); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3040 = i == 8'h31 ? 1'h0 : i == 8'h30 | _GEN_3038; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3042 = i == 8'h32 ? 1'h0 : i == 8'h31 | _GEN_3040; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3043 = i == 8'h59 ? 1'h0 : _GEN_3042; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3044 = i == 8'h5b ? 1'h0 : _GEN_3043; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3045 = i == 8'h62 ? 1'h0 : _GEN_3044; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3047 = i == 8'h65 ? 1'h0 : i == 8'h65 | _GEN_3045; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3048 = i == 8'hb4 ? 1'h0 : _GEN_3047; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3051 = i == 8'hb7 ? 1'h0 : i == 8'hb7 | (i == 8'hb4 | _GEN_3048); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3054 = i == 8'h1 ? 1'h0 : _GEN_2846; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3055 = i == 8'h2 ? 1'h0 : _GEN_3054; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3056 = i == 8'h4 ? 1'h0 : _GEN_3055; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3057 = i == 8'h5 ? 1'h0 : _GEN_3056; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3058 = i == 8'h15 ? 1'h0 : _GEN_3057; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3059 = i == 8'h16 ? 1'h0 : _GEN_3058; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3060 = i == 8'h17 ? 1'h0 : _GEN_3059; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3062 = i == 8'h30 ? 1'h0 : i == 8'h2d | _GEN_3060; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3064 = i == 8'h5a ? 1'h0 : i == 8'h59 | _GEN_3062; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3066 = i == 8'h5b ? 1'h0 : i == 8'h5a | _GEN_3064; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3068 = i == 8'h63 ? 1'h0 : i == 8'h62 | _GEN_3066; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3070 = i == 8'h65 ? 1'h0 : i == 8'h64 | _GEN_3068; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3072 = i == 8'h66 ? 1'h0 : i == 8'h65 | _GEN_3070; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3074 = i == 8'hb4 ? 1'h0 : i == 8'hb4 | _GEN_3072; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3076 = i == 8'hb7 ? 1'h0 : i == 8'hb7 | _GEN_3074; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3077 = i == 8'hc5 ? 1'h0 : _GEN_3076; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3080 = i == 8'hc7 ? 1'h0 : i == 8'hc7 | (i == 8'hc5 | _GEN_3077); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3082 = i == 8'hca ? 1'h0 : i == 8'hca | _GEN_3080; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3085 = i == 8'h1 ? 1'h0 : _GEN_2886; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3086 = i == 8'h2 ? 1'h0 : _GEN_3085; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3087 = i == 8'h4 ? 1'h0 : _GEN_3086; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3088 = i == 8'h5 ? 1'h0 : _GEN_3087; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3089 = i == 8'h16 ? 1'h0 : _GEN_3088; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3090 = i == 8'h17 ? 1'h0 : _GEN_3089; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3091 = i == 8'h2b ? 1'h0 : _GEN_3090; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3092 = i == 8'h30 ? 1'h0 : _GEN_3091; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3093 = i == 8'h58 ? 1'h0 : _GEN_3092; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3096 = i == 8'h5a ? 1'h0 : i == 8'h5a | (i == 8'h58 | _GEN_3093); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3097 = i == 8'h5c ? 1'h0 : _GEN_3096; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3099 = i == 8'h63 ? 1'h0 : i == 8'h5c | _GEN_3097; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3101 = i == 8'hb3 ? 1'h0 : i == 8'h65 | _GEN_3099; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3104 = i == 8'hb4 ? 1'h0 : i == 8'hb4 | (i == 8'hb3 | _GEN_3101); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3106 = i == 8'hb7 ? 1'h0 : i == 8'hb7 | _GEN_3104; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3107 = i == 8'hb8 ? 1'h0 : _GEN_3106; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3109 = i == 8'hc5 ? 1'h0 : i == 8'hb8 | _GEN_3107; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3112 = i == 8'hc6 ? 1'h0 : i == 8'hc6 | (i == 8'hc5 | _GEN_3109); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3113 = i == 8'hc7 ? 1'h0 : _GEN_3112; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3116 = i == 8'hc9 ? 1'h0 : i == 8'hc9 | (i == 8'hc7 | _GEN_3113); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3117 = i == 8'hca ? 1'h0 : _GEN_3116; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3120 = i == 8'hcb ? 1'h0 : i == 8'hcb | (i == 8'hca | _GEN_3117); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3121 = i == 8'hcd ? 1'h0 : _GEN_3120; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3125 = i == 8'h1 ? 1'h0 : i == 8'hba | _GEN_2928; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3126 = i == 8'h2 ? 1'h0 : _GEN_3125; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3127 = i == 8'h4 ? 1'h0 : _GEN_3126; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3128 = i == 8'h5 ? 1'h0 : _GEN_3127; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3131 = i == 8'h2b ? 1'h0 : i == 8'h17 | (i == 8'h16 | _GEN_3128); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3134 = i == 8'h63 ? 1'h0 : i == 8'h62 | (i == 8'h30 | _GEN_3131); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3136 = i == 8'h65 ? 1'h0 : i == 8'h64 | _GEN_3134; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3138 = i == 8'hb1 ? 1'h0 : i == 8'h66 | _GEN_3136; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3140 = i == 8'hb2 ? 1'h0 : i == 8'hb1 | _GEN_3138; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3143 = i == 8'hb3 ? 1'h0 : i == 8'hb3 | (i == 8'hb2 | _GEN_3140); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3145 = i == 8'hb4 ? 1'h0 : i == 8'hb4 | _GEN_3143; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3146 = i == 8'hb5 ? 1'h0 : _GEN_3145; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3148 = i == 8'hb6 ? 1'h0 : i == 8'hb5 | _GEN_3146; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3151 = i == 8'hb7 ? 1'h0 : i == 8'hb7 | (i == 8'hb6 | _GEN_3148); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3153 = i == 8'hb8 ? 1'h0 : i == 8'hb8 | _GEN_3151; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3154 = i == 8'hb9 ? 1'h0 : _GEN_3153; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3156 = i == 8'hba ? 1'h0 : i == 8'hb9 | _GEN_3154; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3158 = i == 8'hc6 ? 1'h0 : i == 8'hba | _GEN_3156; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3161 = i == 8'hc8 ? 1'h0 : i == 8'hc8 | (i == 8'hc6 | _GEN_3158); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3162 = i == 8'hca ? 1'h0 : _GEN_3161; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3165 = i == 8'hcc ? 1'h0 : i == 8'hcc | (i == 8'hca | _GEN_3162); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3166 = i == 8'hce ? 1'h0 : _GEN_3165; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3167 = i == 8'hce | _GEN_3166; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3168 = i == 8'h1 ? 1'h0 : _GEN_2967; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3169 = i == 8'h2 ? 1'h0 : _GEN_3168; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3170 = i == 8'h4 ? 1'h0 : _GEN_3169; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3171 = i == 8'h5 ? 1'h0 : _GEN_3170; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3172 = i == 8'h16 ? 1'h0 : _GEN_3171; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3173 = i == 8'h17 ? 1'h0 : _GEN_3172; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3174 = i == 8'h2b ? 1'h0 : _GEN_3173; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3175 = i == 8'h30 ? 1'h0 : _GEN_3174; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3176 = i == 8'h58 ? 1'h0 : _GEN_3175; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3178 = i == 8'h59 ? 1'h0 : i == 8'h58 | _GEN_3176; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3180 = i == 8'h5a ? 1'h0 : i == 8'h59 | _GEN_3178; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3182 = i == 8'h5b ? 1'h0 : i == 8'h5a | _GEN_3180; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3184 = i == 8'h5c ? 1'h0 : i == 8'h5b | _GEN_3182; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3186 = i == 8'hc5 ? 1'h0 : i == 8'h5c | _GEN_3184; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3189 = i == 8'hc6 ? 1'h0 : i == 8'hc6 | (i == 8'hc5 | _GEN_3186); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3190 = i == 8'hc7 ? 1'h0 : _GEN_3189; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3193 = i == 8'hc8 ? 1'h0 : i == 8'hc8 | (i == 8'hc7 | _GEN_3190); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3194 = i == 8'hc9 ? 1'h0 : _GEN_3193; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3197 = i == 8'hca ? 1'h0 : i == 8'hca | (i == 8'hc9 | _GEN_3194); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3198 = i == 8'hcb ? 1'h0 : _GEN_3197; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3201 = i == 8'hcc ? 1'h0 : i == 8'hcc | (i == 8'hcb | _GEN_3198); // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3202 = i == 8'hcd ? 1'h0 : _GEN_3201; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3206 = i == 8'h1 ? 1'h0 : i == 8'hba | _GEN_3014; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3207 = i == 8'h2 ? 1'h0 : _GEN_3206; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3208 = i == 8'h4 ? 1'h0 : _GEN_3207; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3209 = i == 8'h5 ? 1'h0 : _GEN_3208; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3210 = i == 8'h16 ? 1'h0 : _GEN_3209; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3211 = i == 8'h17 ? 1'h0 : _GEN_3210; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3212 = i == 8'h2b ? 1'h0 : _GEN_3211; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3213 = i == 8'h30 ? 1'h0 : _GEN_3212; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3214 = i == 8'hb1 ? 1'h0 : _GEN_3213; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3216 = i == 8'hb2 ? 1'h0 : i == 8'hb1 | _GEN_3214; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3218 = i == 8'hb3 ? 1'h0 : i == 8'hb2 | _GEN_3216; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3220 = i == 8'hb4 ? 1'h0 : i == 8'hb3 | _GEN_3218; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3222 = i == 8'hb5 ? 1'h0 : i == 8'hb4 | _GEN_3220; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3224 = i == 8'hb6 ? 1'h0 : i == 8'hb5 | _GEN_3222; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3226 = i == 8'hb7 ? 1'h0 : i == 8'hb6 | _GEN_3224; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3228 = i == 8'hb8 ? 1'h0 : i == 8'hb7 | _GEN_3226; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3230 = i == 8'hb9 ? 1'h0 : i == 8'hb8 | _GEN_3228; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3232 = i == 8'hba ? 1'h0 : i == 8'hb9 | _GEN_3230; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3234 = i == 8'hc5 ? 1'h0 : i == 8'hba | _GEN_3232; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3236 = i == 8'hc6 ? 1'h0 : i == 8'hc5 | _GEN_3234; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3238 = i == 8'hc7 ? 1'h0 : i == 8'hc6 | _GEN_3236; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3240 = i == 8'hc8 ? 1'h0 : i == 8'hc7 | _GEN_3238; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3242 = i == 8'hc9 ? 1'h0 : i == 8'hc8 | _GEN_3240; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3244 = i == 8'hca ? 1'h0 : i == 8'hc9 | _GEN_3242; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3246 = i == 8'hcb ? 1'h0 : i == 8'hca | _GEN_3244; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3248 = i == 8'hcc ? 1'h0 : i == 8'hcb | _GEN_3246; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3250 = i == 8'hcd ? 1'h0 : i == 8'hcc | _GEN_3248; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3252 = i == 8'hce ? 1'h0 : i == 8'hcd | _GEN_3250; // @[lut_mem_online.scala 235:34 239:30]
  wire  _GEN_3253 = i == 8'hce | _GEN_3252; // @[lut_mem_online.scala 235:34 239:30]
  wire  _T_3257 = counter < 5'h11; // @[lut_mem_online.scala 250:22]
  wire  _T_3258 = counter < 5'ha; // @[lut_mem_online.scala 255:24]
  wire  _T_3259 = counter >= 5'ha; // @[lut_mem_online.scala 258:30]
  wire [4:0] _outResult_T_1 = counter - 5'ha; // @[lut_mem_online.scala 260:41]
  wire  _GEN_3262 = 3'h1 == _outResult_T_1[2:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_3263 = 3'h2 == _outResult_T_1[2:0] ? buffer_2 : _GEN_3262; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_3264 = 3'h3 == _outResult_T_1[2:0] ? buffer_3 : _GEN_3263; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_3265 = 3'h4 == _outResult_T_1[2:0] ? buffer_4 : _GEN_3264; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_3266 = 3'h5 == _outResult_T_1[2:0] ? buffer_5 : _GEN_3265; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_3267 = 3'h6 == _outResult_T_1[2:0] ? buffer_6 : _GEN_3266; // @[lut_mem_online.scala 260:{23,23}]
  wire  _GEN_3268 = 3'h7 == _outResult_T_1[2:0] ? 1'h0 : _GEN_3267; // @[lut_mem_online.scala 260:{23,23}]
  wire  _T_3263 = ~reset; // @[lut_mem_online.scala 263:21]
  wire  _GEN_3270 = counter >= 5'ha ? _GEN_3268 : outResult; // @[lut_mem_online.scala 258:42 260:23 215:26]
  wire  _GEN_3272 = counter < 5'ha ? 1'h0 : _GEN_3270; // @[lut_mem_online.scala 255:35 257:23]
  wire  _T_3264 = i < 8'h7f; // @[lut_mem_online.scala 274:18]
  wire [9:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 284:24]
  wire [9:0] _i_T_2 = _i_T + 10'h1; // @[lut_mem_online.scala 284:28]
  wire [9:0] _i_T_5 = _i_T + 10'h2; // @[lut_mem_online.scala 286:28]
  wire [9:0] _GEN_3273 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 285:45 286:17 206:18]
  wire [9:0] _GEN_3274 = ~io_inputBit ? _i_T_2 : _GEN_3273; // @[lut_mem_online.scala 283:39 284:17]
  wire  _T_3269 = i < 8'hff; // @[lut_mem_online.scala 289:24]
  wire [7:0] _GEN_3275 = i < 8'hff ? 8'hff : i; // @[lut_mem_online.scala 289:63 297:15 206:18]
  wire [9:0] _GEN_3276 = i < 8'h7f ? _GEN_3274 : {{2'd0}, _GEN_3275}; // @[lut_mem_online.scala 274:61]
  wire [4:0] _counter_T_1 = counter + 5'h1; // @[lut_mem_online.scala 300:30]
  wire  _GEN_3278 = counter < 5'h11 & _GEN_3272; // @[lut_mem_online.scala 250:52 304:21]
  wire [9:0] _GEN_3279 = counter < 5'h11 ? _GEN_3276 : {{2'd0}, i}; // @[lut_mem_online.scala 206:18 250:52]
  wire  _GEN_3302 = io_start & _GEN_3278; // @[lut_mem_online.scala 220:29 327:15]
  wire [9:0] _GEN_3303 = io_start ? _GEN_3279 : 10'h0; // @[lut_mem_online.scala 220:29 325:7]
  wire [9:0] _GEN_5132 = reset ? 10'h0 : _GEN_3303; // @[lut_mem_online.scala 206:{18,18}]
  wire  _GEN_5133 = io_start & _T_3257; // @[lut_mem_online.scala 263:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 334:16]
  always @(posedge clock) begin
    i <= _GEN_5132[7:0]; // @[lut_mem_online.scala 206:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        buffer_0 <= _GEN_3029;
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hc5) begin // @[lut_mem_online.scala 235:34]
          buffer_1 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_1 <= i == 8'hc5 | _GEN_3051;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hcd) begin // @[lut_mem_online.scala 235:34]
          buffer_2 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_2 <= i == 8'hcd | _GEN_3082;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hce) begin // @[lut_mem_online.scala 235:34]
          buffer_3 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_3 <= i == 8'hce | (i == 8'hcd | _GEN_3121);
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        buffer_4 <= _GEN_3167;
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        if (i == 8'hce) begin // @[lut_mem_online.scala 235:34]
          buffer_5 <= 1'h0; // @[lut_mem_online.scala 239:30]
        end else begin
          buffer_5 <= i == 8'hce | (i == 8'hcd | _GEN_3202);
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h8) begin // @[lut_mem_online.scala 232:36]
        buffer_6 <= _GEN_3253;
      end
    end
    if (reset) begin // @[lut_mem_online.scala 212:24]
      counter <= 5'h0; // @[lut_mem_online.scala 212:24]
    end else if (io_start) begin // @[lut_mem_online.scala 220:29]
      if (counter < 5'h11) begin // @[lut_mem_online.scala 250:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 300:19]
      end
    end else begin
      counter <= 5'h0; // @[lut_mem_online.scala 326:13]
    end
    if (reset) begin // @[lut_mem_online.scala 215:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 215:26]
    end else begin
      outResult <= _GEN_3302;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_3257 & ~_T_3258 & _T_3259 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 263:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5133 & _T_3264 & _T_3263) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 277:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5133 & ~_T_3264 & _T_3269 & _T_3263) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 292:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
