module LutMembershipFunctionOnline2_2(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg  buffer_0; // @[lut_mem_online2.scala 76:19]
  reg  buffer_1; // @[lut_mem_online2.scala 76:19]
  reg  buffer_2; // @[lut_mem_online2.scala 76:19]
  reg  buffer_3; // @[lut_mem_online2.scala 76:19]
  reg  buffer_4; // @[lut_mem_online2.scala 76:19]
  reg  buffer_5; // @[lut_mem_online2.scala 76:19]
  reg  buffer_6; // @[lut_mem_online2.scala 76:19]
  reg  buffer_7; // @[lut_mem_online2.scala 76:19]
  reg  buffer_8; // @[lut_mem_online2.scala 76:19]
  reg  buffer_9; // @[lut_mem_online2.scala 76:19]
  reg [6:0] outputBuffer; // @[lut_mem_online2.scala 77:29]
  reg [3:0] counter; // @[lut_mem_online2.scala 79:24]
  reg [3:0] outputCounter; // @[lut_mem_online2.scala 80:30]
  reg  isPassedDelta; // @[lut_mem_online2.scala 82:30]
  reg  isOutputValid; // @[lut_mem_online2.scala 83:30]
  reg  outResult; // @[lut_mem_online2.scala 86:26]
  wire  _GEN_0 = counter == 4'ha | isPassedDelta; // @[lut_mem_online2.scala 114:35 115:25 82:30]
  wire  _T_3 = counter != 4'ha; // @[lut_mem_online2.scala 121:22]
  wire  _GEN_1 = 4'h0 == counter ? io_inputBit : buffer_0; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_2 = 4'h1 == counter ? io_inputBit : buffer_1; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_3 = 4'h2 == counter ? io_inputBit : buffer_2; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_4 = 4'h3 == counter ? io_inputBit : buffer_3; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_5 = 4'h4 == counter ? io_inputBit : buffer_4; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_6 = 4'h5 == counter ? io_inputBit : buffer_5; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_7 = 4'h6 == counter ? io_inputBit : buffer_6; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_8 = 4'h7 == counter ? io_inputBit : buffer_7; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_9 = 4'h8 == counter ? io_inputBit : buffer_8; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _GEN_10 = 4'h9 == counter ? io_inputBit : buffer_9; // @[lut_mem_online2.scala 123:{27,27} 76:19]
  wire  _T_5 = ~reset; // @[lut_mem_online2.scala 127:19]
  wire [3:0] _counter_T_1 = counter + 4'h1; // @[lut_mem_online2.scala 137:30]
  wire  _GEN_11 = counter != 4'ha ? _GEN_1 : buffer_0; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_12 = counter != 4'ha ? _GEN_2 : buffer_1; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_13 = counter != 4'ha ? _GEN_3 : buffer_2; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_14 = counter != 4'ha ? _GEN_4 : buffer_3; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_15 = counter != 4'ha ? _GEN_5 : buffer_4; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_16 = counter != 4'ha ? _GEN_6 : buffer_5; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_17 = counter != 4'ha ? _GEN_7 : buffer_6; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_18 = counter != 4'ha ? _GEN_8 : buffer_7; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_19 = counter != 4'ha ? _GEN_9 : buffer_8; // @[lut_mem_online2.scala 121:38 76:19]
  wire  _GEN_20 = counter != 4'ha ? _GEN_10 : buffer_9; // @[lut_mem_online2.scala 121:38 76:19]
  wire [9:0] _tempCurrentBuf_T = {buffer_9,buffer_8,buffer_7,buffer_6,buffer_5,buffer_4,buffer_3,buffer_2,buffer_1,
    buffer_0}; // @[lut_mem_online2.scala 145:47]
  wire [7:0] _GEN_1085 = {{4'd0}, _tempCurrentBuf_T[7:4]}; // @[Bitwise.scala 108:31]
  wire [7:0] _tempCurrentBuf_T_5 = _GEN_1085 & 8'hf; // @[Bitwise.scala 108:31]
  wire [7:0] _tempCurrentBuf_T_7 = {_tempCurrentBuf_T[3:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _tempCurrentBuf_T_9 = _tempCurrentBuf_T_7 & 8'hf0; // @[Bitwise.scala 108:80]
  wire [7:0] _tempCurrentBuf_T_10 = _tempCurrentBuf_T_5 | _tempCurrentBuf_T_9; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1086 = {{2'd0}, _tempCurrentBuf_T_10[7:2]}; // @[Bitwise.scala 108:31]
  wire [7:0] _tempCurrentBuf_T_15 = _GEN_1086 & 8'h33; // @[Bitwise.scala 108:31]
  wire [7:0] _tempCurrentBuf_T_17 = {_tempCurrentBuf_T_10[5:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _tempCurrentBuf_T_19 = _tempCurrentBuf_T_17 & 8'hcc; // @[Bitwise.scala 108:80]
  wire [7:0] _tempCurrentBuf_T_20 = _tempCurrentBuf_T_15 | _tempCurrentBuf_T_19; // @[Bitwise.scala 108:39]
  wire [7:0] _GEN_1087 = {{1'd0}, _tempCurrentBuf_T_20[7:1]}; // @[Bitwise.scala 108:31]
  wire [7:0] _tempCurrentBuf_T_25 = _GEN_1087 & 8'h55; // @[Bitwise.scala 108:31]
  wire [7:0] _tempCurrentBuf_T_27 = {_tempCurrentBuf_T_20[6:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [7:0] _tempCurrentBuf_T_29 = _tempCurrentBuf_T_27 & 8'haa; // @[Bitwise.scala 108:80]
  wire [7:0] _tempCurrentBuf_T_30 = _tempCurrentBuf_T_25 | _tempCurrentBuf_T_29; // @[Bitwise.scala 108:39]
  wire [9:0] tempCurrentBuf = {_tempCurrentBuf_T_30,_tempCurrentBuf_T[8],_tempCurrentBuf_T[9]}; // @[Cat.scala 33:92]
  wire [6:0] _GEN_223 = 10'hc9 == tempCurrentBuf ? 7'h1 : 7'h0; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_224 = 10'hca == tempCurrentBuf ? 7'h2 : _GEN_223; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_225 = 10'hcb == tempCurrentBuf ? 7'h3 : _GEN_224; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_226 = 10'hcc == tempCurrentBuf ? 7'h4 : _GEN_225; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_227 = 10'hcd == tempCurrentBuf ? 7'h5 : _GEN_226; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_228 = 10'hce == tempCurrentBuf ? 7'h6 : _GEN_227; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_229 = 10'hcf == tempCurrentBuf ? 7'h7 : _GEN_228; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_230 = 10'hd0 == tempCurrentBuf ? 7'h8 : _GEN_229; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_231 = 10'hd1 == tempCurrentBuf ? 7'h9 : _GEN_230; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_232 = 10'hd2 == tempCurrentBuf ? 7'ha : _GEN_231; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_233 = 10'hd3 == tempCurrentBuf ? 7'hb : _GEN_232; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_234 = 10'hd4 == tempCurrentBuf ? 7'hc : _GEN_233; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_235 = 10'hd5 == tempCurrentBuf ? 7'hd : _GEN_234; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_236 = 10'hd6 == tempCurrentBuf ? 7'he : _GEN_235; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_237 = 10'hd7 == tempCurrentBuf ? 7'hf : _GEN_236; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_238 = 10'hd8 == tempCurrentBuf ? 7'h10 : _GEN_237; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_239 = 10'hd9 == tempCurrentBuf ? 7'h11 : _GEN_238; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_240 = 10'hda == tempCurrentBuf ? 7'h12 : _GEN_239; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_241 = 10'hdb == tempCurrentBuf ? 7'h13 : _GEN_240; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_242 = 10'hdc == tempCurrentBuf ? 7'h14 : _GEN_241; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_243 = 10'hdd == tempCurrentBuf ? 7'h15 : _GEN_242; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_244 = 10'hde == tempCurrentBuf ? 7'h16 : _GEN_243; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_245 = 10'hdf == tempCurrentBuf ? 7'h17 : _GEN_244; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_246 = 10'he0 == tempCurrentBuf ? 7'h18 : _GEN_245; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_247 = 10'he1 == tempCurrentBuf ? 7'h19 : _GEN_246; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_248 = 10'he2 == tempCurrentBuf ? 7'h1a : _GEN_247; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_249 = 10'he3 == tempCurrentBuf ? 7'h1b : _GEN_248; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_250 = 10'he4 == tempCurrentBuf ? 7'h1c : _GEN_249; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_251 = 10'he5 == tempCurrentBuf ? 7'h1d : _GEN_250; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_252 = 10'he6 == tempCurrentBuf ? 7'h1e : _GEN_251; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_253 = 10'he7 == tempCurrentBuf ? 7'h1f : _GEN_252; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_254 = 10'he8 == tempCurrentBuf ? 7'h20 : _GEN_253; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_255 = 10'he9 == tempCurrentBuf ? 7'h21 : _GEN_254; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_256 = 10'hea == tempCurrentBuf ? 7'h22 : _GEN_255; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_257 = 10'heb == tempCurrentBuf ? 7'h23 : _GEN_256; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_258 = 10'hec == tempCurrentBuf ? 7'h24 : _GEN_257; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_259 = 10'hed == tempCurrentBuf ? 7'h25 : _GEN_258; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_260 = 10'hee == tempCurrentBuf ? 7'h26 : _GEN_259; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_261 = 10'hef == tempCurrentBuf ? 7'h27 : _GEN_260; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_262 = 10'hf0 == tempCurrentBuf ? 7'h28 : _GEN_261; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_263 = 10'hf1 == tempCurrentBuf ? 7'h29 : _GEN_262; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_264 = 10'hf2 == tempCurrentBuf ? 7'h2a : _GEN_263; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_265 = 10'hf3 == tempCurrentBuf ? 7'h2b : _GEN_264; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_266 = 10'hf4 == tempCurrentBuf ? 7'h2c : _GEN_265; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_267 = 10'hf5 == tempCurrentBuf ? 7'h2d : _GEN_266; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_268 = 10'hf6 == tempCurrentBuf ? 7'h2e : _GEN_267; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_269 = 10'hf7 == tempCurrentBuf ? 7'h2f : _GEN_268; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_270 = 10'hf8 == tempCurrentBuf ? 7'h30 : _GEN_269; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_271 = 10'hf9 == tempCurrentBuf ? 7'h31 : _GEN_270; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_272 = 10'hfa == tempCurrentBuf ? 7'h32 : _GEN_271; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_273 = 10'hfb == tempCurrentBuf ? 7'h33 : _GEN_272; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_274 = 10'hfc == tempCurrentBuf ? 7'h34 : _GEN_273; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_275 = 10'hfd == tempCurrentBuf ? 7'h35 : _GEN_274; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_276 = 10'hfe == tempCurrentBuf ? 7'h36 : _GEN_275; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_277 = 10'hff == tempCurrentBuf ? 7'h37 : _GEN_276; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_278 = 10'h100 == tempCurrentBuf ? 7'h38 : _GEN_277; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_279 = 10'h101 == tempCurrentBuf ? 7'h39 : _GEN_278; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_280 = 10'h102 == tempCurrentBuf ? 7'h3a : _GEN_279; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_281 = 10'h103 == tempCurrentBuf ? 7'h3b : _GEN_280; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_282 = 10'h104 == tempCurrentBuf ? 7'h3c : _GEN_281; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_283 = 10'h105 == tempCurrentBuf ? 7'h3d : _GEN_282; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_284 = 10'h106 == tempCurrentBuf ? 7'h3e : _GEN_283; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_285 = 10'h107 == tempCurrentBuf ? 7'h3f : _GEN_284; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_286 = 10'h108 == tempCurrentBuf ? 7'h40 : _GEN_285; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_287 = 10'h109 == tempCurrentBuf ? 7'h41 : _GEN_286; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_288 = 10'h10a == tempCurrentBuf ? 7'h42 : _GEN_287; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_289 = 10'h10b == tempCurrentBuf ? 7'h43 : _GEN_288; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_290 = 10'h10c == tempCurrentBuf ? 7'h44 : _GEN_289; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_291 = 10'h10d == tempCurrentBuf ? 7'h45 : _GEN_290; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_292 = 10'h10e == tempCurrentBuf ? 7'h46 : _GEN_291; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_293 = 10'h10f == tempCurrentBuf ? 7'h47 : _GEN_292; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_294 = 10'h110 == tempCurrentBuf ? 7'h48 : _GEN_293; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_295 = 10'h111 == tempCurrentBuf ? 7'h49 : _GEN_294; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_296 = 10'h112 == tempCurrentBuf ? 7'h4a : _GEN_295; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_297 = 10'h113 == tempCurrentBuf ? 7'h4b : _GEN_296; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_298 = 10'h114 == tempCurrentBuf ? 7'h4c : _GEN_297; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_299 = 10'h115 == tempCurrentBuf ? 7'h4d : _GEN_298; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_300 = 10'h116 == tempCurrentBuf ? 7'h4e : _GEN_299; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_301 = 10'h117 == tempCurrentBuf ? 7'h4f : _GEN_300; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_302 = 10'h118 == tempCurrentBuf ? 7'h50 : _GEN_301; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_303 = 10'h119 == tempCurrentBuf ? 7'h51 : _GEN_302; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_304 = 10'h11a == tempCurrentBuf ? 7'h52 : _GEN_303; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_305 = 10'h11b == tempCurrentBuf ? 7'h53 : _GEN_304; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_306 = 10'h11c == tempCurrentBuf ? 7'h54 : _GEN_305; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_307 = 10'h11d == tempCurrentBuf ? 7'h55 : _GEN_306; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_308 = 10'h11e == tempCurrentBuf ? 7'h56 : _GEN_307; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_309 = 10'h11f == tempCurrentBuf ? 7'h57 : _GEN_308; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_310 = 10'h120 == tempCurrentBuf ? 7'h58 : _GEN_309; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_311 = 10'h121 == tempCurrentBuf ? 7'h59 : _GEN_310; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_312 = 10'h122 == tempCurrentBuf ? 7'h5a : _GEN_311; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_313 = 10'h123 == tempCurrentBuf ? 7'h5b : _GEN_312; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_314 = 10'h124 == tempCurrentBuf ? 7'h5c : _GEN_313; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_315 = 10'h125 == tempCurrentBuf ? 7'h5d : _GEN_314; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_316 = 10'h126 == tempCurrentBuf ? 7'h5e : _GEN_315; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_317 = 10'h127 == tempCurrentBuf ? 7'h5f : _GEN_316; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_318 = 10'h128 == tempCurrentBuf ? 7'h60 : _GEN_317; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_319 = 10'h129 == tempCurrentBuf ? 7'h61 : _GEN_318; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_320 = 10'h12a == tempCurrentBuf ? 7'h62 : _GEN_319; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_321 = 10'h12b == tempCurrentBuf ? 7'h63 : _GEN_320; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_322 = 10'h12c == tempCurrentBuf ? 7'h64 : _GEN_321; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_323 = 10'h12d == tempCurrentBuf ? 7'h0 : _GEN_322; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_324 = 10'h12e == tempCurrentBuf ? 7'h0 : _GEN_323; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_325 = 10'h12f == tempCurrentBuf ? 7'h0 : _GEN_324; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_326 = 10'h130 == tempCurrentBuf ? 7'h0 : _GEN_325; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_327 = 10'h131 == tempCurrentBuf ? 7'h0 : _GEN_326; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_328 = 10'h132 == tempCurrentBuf ? 7'h0 : _GEN_327; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_329 = 10'h133 == tempCurrentBuf ? 7'h0 : _GEN_328; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_330 = 10'h134 == tempCurrentBuf ? 7'h0 : _GEN_329; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_331 = 10'h135 == tempCurrentBuf ? 7'h0 : _GEN_330; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_332 = 10'h136 == tempCurrentBuf ? 7'h0 : _GEN_331; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_333 = 10'h137 == tempCurrentBuf ? 7'h0 : _GEN_332; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_334 = 10'h138 == tempCurrentBuf ? 7'h0 : _GEN_333; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_335 = 10'h139 == tempCurrentBuf ? 7'h0 : _GEN_334; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_336 = 10'h13a == tempCurrentBuf ? 7'h0 : _GEN_335; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_337 = 10'h13b == tempCurrentBuf ? 7'h0 : _GEN_336; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_338 = 10'h13c == tempCurrentBuf ? 7'h0 : _GEN_337; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_339 = 10'h13d == tempCurrentBuf ? 7'h0 : _GEN_338; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_340 = 10'h13e == tempCurrentBuf ? 7'h0 : _GEN_339; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_341 = 10'h13f == tempCurrentBuf ? 7'h0 : _GEN_340; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_342 = 10'h140 == tempCurrentBuf ? 7'h0 : _GEN_341; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_343 = 10'h141 == tempCurrentBuf ? 7'h0 : _GEN_342; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_344 = 10'h142 == tempCurrentBuf ? 7'h0 : _GEN_343; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_345 = 10'h143 == tempCurrentBuf ? 7'h0 : _GEN_344; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_346 = 10'h144 == tempCurrentBuf ? 7'h0 : _GEN_345; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_347 = 10'h145 == tempCurrentBuf ? 7'h0 : _GEN_346; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_348 = 10'h146 == tempCurrentBuf ? 7'h0 : _GEN_347; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_349 = 10'h147 == tempCurrentBuf ? 7'h0 : _GEN_348; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_350 = 10'h148 == tempCurrentBuf ? 7'h0 : _GEN_349; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_351 = 10'h149 == tempCurrentBuf ? 7'h0 : _GEN_350; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_352 = 10'h14a == tempCurrentBuf ? 7'h0 : _GEN_351; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_353 = 10'h14b == tempCurrentBuf ? 7'h0 : _GEN_352; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_354 = 10'h14c == tempCurrentBuf ? 7'h0 : _GEN_353; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_355 = 10'h14d == tempCurrentBuf ? 7'h0 : _GEN_354; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_356 = 10'h14e == tempCurrentBuf ? 7'h0 : _GEN_355; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_357 = 10'h14f == tempCurrentBuf ? 7'h0 : _GEN_356; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_358 = 10'h150 == tempCurrentBuf ? 7'h0 : _GEN_357; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_359 = 10'h151 == tempCurrentBuf ? 7'h0 : _GEN_358; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_360 = 10'h152 == tempCurrentBuf ? 7'h0 : _GEN_359; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_361 = 10'h153 == tempCurrentBuf ? 7'h0 : _GEN_360; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_362 = 10'h154 == tempCurrentBuf ? 7'h0 : _GEN_361; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_363 = 10'h155 == tempCurrentBuf ? 7'h0 : _GEN_362; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_364 = 10'h156 == tempCurrentBuf ? 7'h0 : _GEN_363; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_365 = 10'h157 == tempCurrentBuf ? 7'h0 : _GEN_364; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_366 = 10'h158 == tempCurrentBuf ? 7'h0 : _GEN_365; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_367 = 10'h159 == tempCurrentBuf ? 7'h0 : _GEN_366; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_368 = 10'h15a == tempCurrentBuf ? 7'h0 : _GEN_367; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_369 = 10'h15b == tempCurrentBuf ? 7'h0 : _GEN_368; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_370 = 10'h15c == tempCurrentBuf ? 7'h0 : _GEN_369; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_371 = 10'h15d == tempCurrentBuf ? 7'h0 : _GEN_370; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_372 = 10'h15e == tempCurrentBuf ? 7'h0 : _GEN_371; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_373 = 10'h15f == tempCurrentBuf ? 7'h0 : _GEN_372; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_374 = 10'h160 == tempCurrentBuf ? 7'h0 : _GEN_373; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_375 = 10'h161 == tempCurrentBuf ? 7'h0 : _GEN_374; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_376 = 10'h162 == tempCurrentBuf ? 7'h0 : _GEN_375; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_377 = 10'h163 == tempCurrentBuf ? 7'h0 : _GEN_376; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_378 = 10'h164 == tempCurrentBuf ? 7'h0 : _GEN_377; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_379 = 10'h165 == tempCurrentBuf ? 7'h0 : _GEN_378; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_380 = 10'h166 == tempCurrentBuf ? 7'h0 : _GEN_379; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_381 = 10'h167 == tempCurrentBuf ? 7'h0 : _GEN_380; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_382 = 10'h168 == tempCurrentBuf ? 7'h0 : _GEN_381; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_383 = 10'h169 == tempCurrentBuf ? 7'h0 : _GEN_382; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_384 = 10'h16a == tempCurrentBuf ? 7'h0 : _GEN_383; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_385 = 10'h16b == tempCurrentBuf ? 7'h0 : _GEN_384; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_386 = 10'h16c == tempCurrentBuf ? 7'h0 : _GEN_385; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_387 = 10'h16d == tempCurrentBuf ? 7'h0 : _GEN_386; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_388 = 10'h16e == tempCurrentBuf ? 7'h0 : _GEN_387; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_389 = 10'h16f == tempCurrentBuf ? 7'h0 : _GEN_388; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_390 = 10'h170 == tempCurrentBuf ? 7'h0 : _GEN_389; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_391 = 10'h171 == tempCurrentBuf ? 7'h0 : _GEN_390; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_392 = 10'h172 == tempCurrentBuf ? 7'h0 : _GEN_391; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_393 = 10'h173 == tempCurrentBuf ? 7'h0 : _GEN_392; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_394 = 10'h174 == tempCurrentBuf ? 7'h0 : _GEN_393; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_395 = 10'h175 == tempCurrentBuf ? 7'h0 : _GEN_394; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_396 = 10'h176 == tempCurrentBuf ? 7'h0 : _GEN_395; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_397 = 10'h177 == tempCurrentBuf ? 7'h0 : _GEN_396; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_398 = 10'h178 == tempCurrentBuf ? 7'h0 : _GEN_397; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_399 = 10'h179 == tempCurrentBuf ? 7'h0 : _GEN_398; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_400 = 10'h17a == tempCurrentBuf ? 7'h0 : _GEN_399; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_401 = 10'h17b == tempCurrentBuf ? 7'h0 : _GEN_400; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_402 = 10'h17c == tempCurrentBuf ? 7'h0 : _GEN_401; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_403 = 10'h17d == tempCurrentBuf ? 7'h0 : _GEN_402; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_404 = 10'h17e == tempCurrentBuf ? 7'h0 : _GEN_403; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_405 = 10'h17f == tempCurrentBuf ? 7'h0 : _GEN_404; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_406 = 10'h180 == tempCurrentBuf ? 7'h0 : _GEN_405; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_407 = 10'h181 == tempCurrentBuf ? 7'h0 : _GEN_406; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_408 = 10'h182 == tempCurrentBuf ? 7'h0 : _GEN_407; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_409 = 10'h183 == tempCurrentBuf ? 7'h0 : _GEN_408; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_410 = 10'h184 == tempCurrentBuf ? 7'h0 : _GEN_409; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_411 = 10'h185 == tempCurrentBuf ? 7'h0 : _GEN_410; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_412 = 10'h186 == tempCurrentBuf ? 7'h0 : _GEN_411; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_413 = 10'h187 == tempCurrentBuf ? 7'h0 : _GEN_412; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_414 = 10'h188 == tempCurrentBuf ? 7'h0 : _GEN_413; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_415 = 10'h189 == tempCurrentBuf ? 7'h0 : _GEN_414; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_416 = 10'h18a == tempCurrentBuf ? 7'h0 : _GEN_415; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_417 = 10'h18b == tempCurrentBuf ? 7'h0 : _GEN_416; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_418 = 10'h18c == tempCurrentBuf ? 7'h0 : _GEN_417; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_419 = 10'h18d == tempCurrentBuf ? 7'h0 : _GEN_418; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_420 = 10'h18e == tempCurrentBuf ? 7'h0 : _GEN_419; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_421 = 10'h18f == tempCurrentBuf ? 7'h0 : _GEN_420; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_422 = 10'h190 == tempCurrentBuf ? 7'h0 : _GEN_421; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_423 = 10'h191 == tempCurrentBuf ? 7'h0 : _GEN_422; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_424 = 10'h192 == tempCurrentBuf ? 7'h0 : _GEN_423; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_425 = 10'h193 == tempCurrentBuf ? 7'h0 : _GEN_424; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_426 = 10'h194 == tempCurrentBuf ? 7'h0 : _GEN_425; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_427 = 10'h195 == tempCurrentBuf ? 7'h0 : _GEN_426; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_428 = 10'h196 == tempCurrentBuf ? 7'h0 : _GEN_427; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_429 = 10'h197 == tempCurrentBuf ? 7'h0 : _GEN_428; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_430 = 10'h198 == tempCurrentBuf ? 7'h0 : _GEN_429; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_431 = 10'h199 == tempCurrentBuf ? 7'h0 : _GEN_430; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_432 = 10'h19a == tempCurrentBuf ? 7'h0 : _GEN_431; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_433 = 10'h19b == tempCurrentBuf ? 7'h0 : _GEN_432; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_434 = 10'h19c == tempCurrentBuf ? 7'h0 : _GEN_433; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_435 = 10'h19d == tempCurrentBuf ? 7'h0 : _GEN_434; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_436 = 10'h19e == tempCurrentBuf ? 7'h0 : _GEN_435; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_437 = 10'h19f == tempCurrentBuf ? 7'h0 : _GEN_436; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_438 = 10'h1a0 == tempCurrentBuf ? 7'h0 : _GEN_437; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_439 = 10'h1a1 == tempCurrentBuf ? 7'h0 : _GEN_438; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_440 = 10'h1a2 == tempCurrentBuf ? 7'h0 : _GEN_439; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_441 = 10'h1a3 == tempCurrentBuf ? 7'h0 : _GEN_440; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_442 = 10'h1a4 == tempCurrentBuf ? 7'h0 : _GEN_441; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_443 = 10'h1a5 == tempCurrentBuf ? 7'h0 : _GEN_442; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_444 = 10'h1a6 == tempCurrentBuf ? 7'h0 : _GEN_443; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_445 = 10'h1a7 == tempCurrentBuf ? 7'h0 : _GEN_444; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_446 = 10'h1a8 == tempCurrentBuf ? 7'h0 : _GEN_445; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_447 = 10'h1a9 == tempCurrentBuf ? 7'h0 : _GEN_446; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_448 = 10'h1aa == tempCurrentBuf ? 7'h0 : _GEN_447; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_449 = 10'h1ab == tempCurrentBuf ? 7'h0 : _GEN_448; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_450 = 10'h1ac == tempCurrentBuf ? 7'h0 : _GEN_449; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_451 = 10'h1ad == tempCurrentBuf ? 7'h0 : _GEN_450; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_452 = 10'h1ae == tempCurrentBuf ? 7'h0 : _GEN_451; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_453 = 10'h1af == tempCurrentBuf ? 7'h0 : _GEN_452; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_454 = 10'h1b0 == tempCurrentBuf ? 7'h0 : _GEN_453; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_455 = 10'h1b1 == tempCurrentBuf ? 7'h0 : _GEN_454; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_456 = 10'h1b2 == tempCurrentBuf ? 7'h0 : _GEN_455; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_457 = 10'h1b3 == tempCurrentBuf ? 7'h0 : _GEN_456; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_458 = 10'h1b4 == tempCurrentBuf ? 7'h0 : _GEN_457; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_459 = 10'h1b5 == tempCurrentBuf ? 7'h0 : _GEN_458; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_460 = 10'h1b6 == tempCurrentBuf ? 7'h0 : _GEN_459; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_461 = 10'h1b7 == tempCurrentBuf ? 7'h0 : _GEN_460; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_462 = 10'h1b8 == tempCurrentBuf ? 7'h0 : _GEN_461; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_463 = 10'h1b9 == tempCurrentBuf ? 7'h0 : _GEN_462; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_464 = 10'h1ba == tempCurrentBuf ? 7'h0 : _GEN_463; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_465 = 10'h1bb == tempCurrentBuf ? 7'h0 : _GEN_464; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_466 = 10'h1bc == tempCurrentBuf ? 7'h0 : _GEN_465; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_467 = 10'h1bd == tempCurrentBuf ? 7'h0 : _GEN_466; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_468 = 10'h1be == tempCurrentBuf ? 7'h0 : _GEN_467; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_469 = 10'h1bf == tempCurrentBuf ? 7'h0 : _GEN_468; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_470 = 10'h1c0 == tempCurrentBuf ? 7'h0 : _GEN_469; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_471 = 10'h1c1 == tempCurrentBuf ? 7'h0 : _GEN_470; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_472 = 10'h1c2 == tempCurrentBuf ? 7'h0 : _GEN_471; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_473 = 10'h1c3 == tempCurrentBuf ? 7'h0 : _GEN_472; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_474 = 10'h1c4 == tempCurrentBuf ? 7'h0 : _GEN_473; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_475 = 10'h1c5 == tempCurrentBuf ? 7'h0 : _GEN_474; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_476 = 10'h1c6 == tempCurrentBuf ? 7'h0 : _GEN_475; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_477 = 10'h1c7 == tempCurrentBuf ? 7'h0 : _GEN_476; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_478 = 10'h1c8 == tempCurrentBuf ? 7'h0 : _GEN_477; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_479 = 10'h1c9 == tempCurrentBuf ? 7'h0 : _GEN_478; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_480 = 10'h1ca == tempCurrentBuf ? 7'h0 : _GEN_479; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_481 = 10'h1cb == tempCurrentBuf ? 7'h0 : _GEN_480; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_482 = 10'h1cc == tempCurrentBuf ? 7'h0 : _GEN_481; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_483 = 10'h1cd == tempCurrentBuf ? 7'h0 : _GEN_482; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_484 = 10'h1ce == tempCurrentBuf ? 7'h0 : _GEN_483; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_485 = 10'h1cf == tempCurrentBuf ? 7'h0 : _GEN_484; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_486 = 10'h1d0 == tempCurrentBuf ? 7'h0 : _GEN_485; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_487 = 10'h1d1 == tempCurrentBuf ? 7'h0 : _GEN_486; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_488 = 10'h1d2 == tempCurrentBuf ? 7'h0 : _GEN_487; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_489 = 10'h1d3 == tempCurrentBuf ? 7'h0 : _GEN_488; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_490 = 10'h1d4 == tempCurrentBuf ? 7'h0 : _GEN_489; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_491 = 10'h1d5 == tempCurrentBuf ? 7'h0 : _GEN_490; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_492 = 10'h1d6 == tempCurrentBuf ? 7'h0 : _GEN_491; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_493 = 10'h1d7 == tempCurrentBuf ? 7'h0 : _GEN_492; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_494 = 10'h1d8 == tempCurrentBuf ? 7'h0 : _GEN_493; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_495 = 10'h1d9 == tempCurrentBuf ? 7'h0 : _GEN_494; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_496 = 10'h1da == tempCurrentBuf ? 7'h0 : _GEN_495; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_497 = 10'h1db == tempCurrentBuf ? 7'h0 : _GEN_496; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_498 = 10'h1dc == tempCurrentBuf ? 7'h0 : _GEN_497; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_499 = 10'h1dd == tempCurrentBuf ? 7'h0 : _GEN_498; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_500 = 10'h1de == tempCurrentBuf ? 7'h0 : _GEN_499; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_501 = 10'h1df == tempCurrentBuf ? 7'h0 : _GEN_500; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_502 = 10'h1e0 == tempCurrentBuf ? 7'h0 : _GEN_501; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_503 = 10'h1e1 == tempCurrentBuf ? 7'h0 : _GEN_502; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_504 = 10'h1e2 == tempCurrentBuf ? 7'h0 : _GEN_503; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_505 = 10'h1e3 == tempCurrentBuf ? 7'h0 : _GEN_504; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_506 = 10'h1e4 == tempCurrentBuf ? 7'h0 : _GEN_505; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_507 = 10'h1e5 == tempCurrentBuf ? 7'h0 : _GEN_506; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_508 = 10'h1e6 == tempCurrentBuf ? 7'h0 : _GEN_507; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_509 = 10'h1e7 == tempCurrentBuf ? 7'h0 : _GEN_508; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_510 = 10'h1e8 == tempCurrentBuf ? 7'h0 : _GEN_509; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_511 = 10'h1e9 == tempCurrentBuf ? 7'h0 : _GEN_510; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_512 = 10'h1ea == tempCurrentBuf ? 7'h0 : _GEN_511; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_513 = 10'h1eb == tempCurrentBuf ? 7'h0 : _GEN_512; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_514 = 10'h1ec == tempCurrentBuf ? 7'h0 : _GEN_513; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_515 = 10'h1ed == tempCurrentBuf ? 7'h0 : _GEN_514; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_516 = 10'h1ee == tempCurrentBuf ? 7'h0 : _GEN_515; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_517 = 10'h1ef == tempCurrentBuf ? 7'h0 : _GEN_516; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_518 = 10'h1f0 == tempCurrentBuf ? 7'h0 : _GEN_517; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_519 = 10'h1f1 == tempCurrentBuf ? 7'h0 : _GEN_518; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_520 = 10'h1f2 == tempCurrentBuf ? 7'h0 : _GEN_519; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_521 = 10'h1f3 == tempCurrentBuf ? 7'h0 : _GEN_520; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_522 = 10'h1f4 == tempCurrentBuf ? 7'h0 : _GEN_521; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_523 = 10'h1f5 == tempCurrentBuf ? 7'h0 : _GEN_522; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_524 = 10'h1f6 == tempCurrentBuf ? 7'h0 : _GEN_523; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_525 = 10'h1f7 == tempCurrentBuf ? 7'h0 : _GEN_524; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_526 = 10'h1f8 == tempCurrentBuf ? 7'h0 : _GEN_525; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_527 = 10'h1f9 == tempCurrentBuf ? 7'h0 : _GEN_526; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_528 = 10'h1fa == tempCurrentBuf ? 7'h0 : _GEN_527; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_529 = 10'h1fb == tempCurrentBuf ? 7'h0 : _GEN_528; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_530 = 10'h1fc == tempCurrentBuf ? 7'h0 : _GEN_529; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_531 = 10'h1fd == tempCurrentBuf ? 7'h0 : _GEN_530; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_532 = 10'h1fe == tempCurrentBuf ? 7'h0 : _GEN_531; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_533 = 10'h1ff == tempCurrentBuf ? 7'h0 : _GEN_532; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_534 = 10'h200 == tempCurrentBuf ? 7'h0 : _GEN_533; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_535 = 10'h201 == tempCurrentBuf ? 7'h0 : _GEN_534; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_536 = 10'h202 == tempCurrentBuf ? 7'h0 : _GEN_535; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_537 = 10'h203 == tempCurrentBuf ? 7'h0 : _GEN_536; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_538 = 10'h204 == tempCurrentBuf ? 7'h0 : _GEN_537; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_539 = 10'h205 == tempCurrentBuf ? 7'h0 : _GEN_538; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_540 = 10'h206 == tempCurrentBuf ? 7'h0 : _GEN_539; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_541 = 10'h207 == tempCurrentBuf ? 7'h0 : _GEN_540; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_542 = 10'h208 == tempCurrentBuf ? 7'h0 : _GEN_541; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_543 = 10'h209 == tempCurrentBuf ? 7'h0 : _GEN_542; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_544 = 10'h20a == tempCurrentBuf ? 7'h0 : _GEN_543; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_545 = 10'h20b == tempCurrentBuf ? 7'h0 : _GEN_544; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_546 = 10'h20c == tempCurrentBuf ? 7'h0 : _GEN_545; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_547 = 10'h20d == tempCurrentBuf ? 7'h0 : _GEN_546; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_548 = 10'h20e == tempCurrentBuf ? 7'h0 : _GEN_547; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_549 = 10'h20f == tempCurrentBuf ? 7'h0 : _GEN_548; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_550 = 10'h210 == tempCurrentBuf ? 7'h0 : _GEN_549; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_551 = 10'h211 == tempCurrentBuf ? 7'h0 : _GEN_550; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_552 = 10'h212 == tempCurrentBuf ? 7'h0 : _GEN_551; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_553 = 10'h213 == tempCurrentBuf ? 7'h0 : _GEN_552; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_554 = 10'h214 == tempCurrentBuf ? 7'h0 : _GEN_553; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_555 = 10'h215 == tempCurrentBuf ? 7'h0 : _GEN_554; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_556 = 10'h216 == tempCurrentBuf ? 7'h0 : _GEN_555; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_557 = 10'h217 == tempCurrentBuf ? 7'h0 : _GEN_556; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_558 = 10'h218 == tempCurrentBuf ? 7'h0 : _GEN_557; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_559 = 10'h219 == tempCurrentBuf ? 7'h0 : _GEN_558; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_560 = 10'h21a == tempCurrentBuf ? 7'h0 : _GEN_559; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_561 = 10'h21b == tempCurrentBuf ? 7'h0 : _GEN_560; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_562 = 10'h21c == tempCurrentBuf ? 7'h0 : _GEN_561; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_563 = 10'h21d == tempCurrentBuf ? 7'h0 : _GEN_562; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_564 = 10'h21e == tempCurrentBuf ? 7'h0 : _GEN_563; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_565 = 10'h21f == tempCurrentBuf ? 7'h0 : _GEN_564; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_566 = 10'h220 == tempCurrentBuf ? 7'h0 : _GEN_565; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_567 = 10'h221 == tempCurrentBuf ? 7'h0 : _GEN_566; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_568 = 10'h222 == tempCurrentBuf ? 7'h0 : _GEN_567; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_569 = 10'h223 == tempCurrentBuf ? 7'h0 : _GEN_568; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_570 = 10'h224 == tempCurrentBuf ? 7'h0 : _GEN_569; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_571 = 10'h225 == tempCurrentBuf ? 7'h0 : _GEN_570; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_572 = 10'h226 == tempCurrentBuf ? 7'h0 : _GEN_571; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_573 = 10'h227 == tempCurrentBuf ? 7'h0 : _GEN_572; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_574 = 10'h228 == tempCurrentBuf ? 7'h0 : _GEN_573; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_575 = 10'h229 == tempCurrentBuf ? 7'h0 : _GEN_574; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_576 = 10'h22a == tempCurrentBuf ? 7'h0 : _GEN_575; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_577 = 10'h22b == tempCurrentBuf ? 7'h0 : _GEN_576; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_578 = 10'h22c == tempCurrentBuf ? 7'h0 : _GEN_577; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_579 = 10'h22d == tempCurrentBuf ? 7'h0 : _GEN_578; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_580 = 10'h22e == tempCurrentBuf ? 7'h0 : _GEN_579; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_581 = 10'h22f == tempCurrentBuf ? 7'h0 : _GEN_580; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_582 = 10'h230 == tempCurrentBuf ? 7'h0 : _GEN_581; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_583 = 10'h231 == tempCurrentBuf ? 7'h0 : _GEN_582; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_584 = 10'h232 == tempCurrentBuf ? 7'h0 : _GEN_583; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_585 = 10'h233 == tempCurrentBuf ? 7'h0 : _GEN_584; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_586 = 10'h234 == tempCurrentBuf ? 7'h0 : _GEN_585; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_587 = 10'h235 == tempCurrentBuf ? 7'h0 : _GEN_586; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_588 = 10'h236 == tempCurrentBuf ? 7'h0 : _GEN_587; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_589 = 10'h237 == tempCurrentBuf ? 7'h0 : _GEN_588; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_590 = 10'h238 == tempCurrentBuf ? 7'h0 : _GEN_589; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_591 = 10'h239 == tempCurrentBuf ? 7'h0 : _GEN_590; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_592 = 10'h23a == tempCurrentBuf ? 7'h0 : _GEN_591; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_593 = 10'h23b == tempCurrentBuf ? 7'h0 : _GEN_592; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_594 = 10'h23c == tempCurrentBuf ? 7'h0 : _GEN_593; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_595 = 10'h23d == tempCurrentBuf ? 7'h0 : _GEN_594; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_596 = 10'h23e == tempCurrentBuf ? 7'h0 : _GEN_595; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_597 = 10'h23f == tempCurrentBuf ? 7'h0 : _GEN_596; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_598 = 10'h240 == tempCurrentBuf ? 7'h0 : _GEN_597; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_599 = 10'h241 == tempCurrentBuf ? 7'h0 : _GEN_598; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_600 = 10'h242 == tempCurrentBuf ? 7'h0 : _GEN_599; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_601 = 10'h243 == tempCurrentBuf ? 7'h0 : _GEN_600; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_602 = 10'h244 == tempCurrentBuf ? 7'h0 : _GEN_601; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_603 = 10'h245 == tempCurrentBuf ? 7'h0 : _GEN_602; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_604 = 10'h246 == tempCurrentBuf ? 7'h0 : _GEN_603; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_605 = 10'h247 == tempCurrentBuf ? 7'h0 : _GEN_604; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_606 = 10'h248 == tempCurrentBuf ? 7'h0 : _GEN_605; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_607 = 10'h249 == tempCurrentBuf ? 7'h0 : _GEN_606; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_608 = 10'h24a == tempCurrentBuf ? 7'h0 : _GEN_607; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_609 = 10'h24b == tempCurrentBuf ? 7'h0 : _GEN_608; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_610 = 10'h24c == tempCurrentBuf ? 7'h0 : _GEN_609; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_611 = 10'h24d == tempCurrentBuf ? 7'h0 : _GEN_610; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_612 = 10'h24e == tempCurrentBuf ? 7'h0 : _GEN_611; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_613 = 10'h24f == tempCurrentBuf ? 7'h0 : _GEN_612; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_614 = 10'h250 == tempCurrentBuf ? 7'h0 : _GEN_613; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_615 = 10'h251 == tempCurrentBuf ? 7'h0 : _GEN_614; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_616 = 10'h252 == tempCurrentBuf ? 7'h0 : _GEN_615; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_617 = 10'h253 == tempCurrentBuf ? 7'h0 : _GEN_616; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_618 = 10'h254 == tempCurrentBuf ? 7'h0 : _GEN_617; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_619 = 10'h255 == tempCurrentBuf ? 7'h0 : _GEN_618; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_620 = 10'h256 == tempCurrentBuf ? 7'h0 : _GEN_619; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_621 = 10'h257 == tempCurrentBuf ? 7'h0 : _GEN_620; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_622 = 10'h258 == tempCurrentBuf ? 7'h0 : _GEN_621; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_623 = 10'h259 == tempCurrentBuf ? 7'h0 : _GEN_622; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_624 = 10'h25a == tempCurrentBuf ? 7'h0 : _GEN_623; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_625 = 10'h25b == tempCurrentBuf ? 7'h0 : _GEN_624; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_626 = 10'h25c == tempCurrentBuf ? 7'h0 : _GEN_625; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_627 = 10'h25d == tempCurrentBuf ? 7'h0 : _GEN_626; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_628 = 10'h25e == tempCurrentBuf ? 7'h0 : _GEN_627; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_629 = 10'h25f == tempCurrentBuf ? 7'h0 : _GEN_628; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_630 = 10'h260 == tempCurrentBuf ? 7'h0 : _GEN_629; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_631 = 10'h261 == tempCurrentBuf ? 7'h0 : _GEN_630; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_632 = 10'h262 == tempCurrentBuf ? 7'h0 : _GEN_631; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_633 = 10'h263 == tempCurrentBuf ? 7'h0 : _GEN_632; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_634 = 10'h264 == tempCurrentBuf ? 7'h0 : _GEN_633; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_635 = 10'h265 == tempCurrentBuf ? 7'h0 : _GEN_634; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_636 = 10'h266 == tempCurrentBuf ? 7'h0 : _GEN_635; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_637 = 10'h267 == tempCurrentBuf ? 7'h0 : _GEN_636; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_638 = 10'h268 == tempCurrentBuf ? 7'h0 : _GEN_637; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_639 = 10'h269 == tempCurrentBuf ? 7'h0 : _GEN_638; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_640 = 10'h26a == tempCurrentBuf ? 7'h0 : _GEN_639; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_641 = 10'h26b == tempCurrentBuf ? 7'h0 : _GEN_640; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_642 = 10'h26c == tempCurrentBuf ? 7'h0 : _GEN_641; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_643 = 10'h26d == tempCurrentBuf ? 7'h0 : _GEN_642; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_644 = 10'h26e == tempCurrentBuf ? 7'h0 : _GEN_643; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_645 = 10'h26f == tempCurrentBuf ? 7'h0 : _GEN_644; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_646 = 10'h270 == tempCurrentBuf ? 7'h0 : _GEN_645; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_647 = 10'h271 == tempCurrentBuf ? 7'h0 : _GEN_646; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_648 = 10'h272 == tempCurrentBuf ? 7'h0 : _GEN_647; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_649 = 10'h273 == tempCurrentBuf ? 7'h0 : _GEN_648; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_650 = 10'h274 == tempCurrentBuf ? 7'h0 : _GEN_649; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_651 = 10'h275 == tempCurrentBuf ? 7'h0 : _GEN_650; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_652 = 10'h276 == tempCurrentBuf ? 7'h0 : _GEN_651; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_653 = 10'h277 == tempCurrentBuf ? 7'h0 : _GEN_652; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_654 = 10'h278 == tempCurrentBuf ? 7'h0 : _GEN_653; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_655 = 10'h279 == tempCurrentBuf ? 7'h0 : _GEN_654; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_656 = 10'h27a == tempCurrentBuf ? 7'h0 : _GEN_655; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_657 = 10'h27b == tempCurrentBuf ? 7'h0 : _GEN_656; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_658 = 10'h27c == tempCurrentBuf ? 7'h0 : _GEN_657; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_659 = 10'h27d == tempCurrentBuf ? 7'h0 : _GEN_658; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_660 = 10'h27e == tempCurrentBuf ? 7'h0 : _GEN_659; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_661 = 10'h27f == tempCurrentBuf ? 7'h0 : _GEN_660; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_662 = 10'h280 == tempCurrentBuf ? 7'h0 : _GEN_661; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_663 = 10'h281 == tempCurrentBuf ? 7'h0 : _GEN_662; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_664 = 10'h282 == tempCurrentBuf ? 7'h0 : _GEN_663; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_665 = 10'h283 == tempCurrentBuf ? 7'h0 : _GEN_664; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_666 = 10'h284 == tempCurrentBuf ? 7'h0 : _GEN_665; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_667 = 10'h285 == tempCurrentBuf ? 7'h0 : _GEN_666; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_668 = 10'h286 == tempCurrentBuf ? 7'h0 : _GEN_667; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_669 = 10'h287 == tempCurrentBuf ? 7'h0 : _GEN_668; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_670 = 10'h288 == tempCurrentBuf ? 7'h0 : _GEN_669; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_671 = 10'h289 == tempCurrentBuf ? 7'h0 : _GEN_670; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_672 = 10'h28a == tempCurrentBuf ? 7'h0 : _GEN_671; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_673 = 10'h28b == tempCurrentBuf ? 7'h0 : _GEN_672; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_674 = 10'h28c == tempCurrentBuf ? 7'h0 : _GEN_673; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_675 = 10'h28d == tempCurrentBuf ? 7'h0 : _GEN_674; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_676 = 10'h28e == tempCurrentBuf ? 7'h0 : _GEN_675; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_677 = 10'h28f == tempCurrentBuf ? 7'h0 : _GEN_676; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_678 = 10'h290 == tempCurrentBuf ? 7'h0 : _GEN_677; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_679 = 10'h291 == tempCurrentBuf ? 7'h0 : _GEN_678; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_680 = 10'h292 == tempCurrentBuf ? 7'h0 : _GEN_679; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_681 = 10'h293 == tempCurrentBuf ? 7'h0 : _GEN_680; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_682 = 10'h294 == tempCurrentBuf ? 7'h0 : _GEN_681; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_683 = 10'h295 == tempCurrentBuf ? 7'h0 : _GEN_682; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_684 = 10'h296 == tempCurrentBuf ? 7'h0 : _GEN_683; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_685 = 10'h297 == tempCurrentBuf ? 7'h0 : _GEN_684; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_686 = 10'h298 == tempCurrentBuf ? 7'h0 : _GEN_685; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_687 = 10'h299 == tempCurrentBuf ? 7'h0 : _GEN_686; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_688 = 10'h29a == tempCurrentBuf ? 7'h0 : _GEN_687; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_689 = 10'h29b == tempCurrentBuf ? 7'h0 : _GEN_688; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_690 = 10'h29c == tempCurrentBuf ? 7'h0 : _GEN_689; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_691 = 10'h29d == tempCurrentBuf ? 7'h0 : _GEN_690; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_692 = 10'h29e == tempCurrentBuf ? 7'h0 : _GEN_691; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_693 = 10'h29f == tempCurrentBuf ? 7'h0 : _GEN_692; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_694 = 10'h2a0 == tempCurrentBuf ? 7'h0 : _GEN_693; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_695 = 10'h2a1 == tempCurrentBuf ? 7'h0 : _GEN_694; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_696 = 10'h2a2 == tempCurrentBuf ? 7'h0 : _GEN_695; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_697 = 10'h2a3 == tempCurrentBuf ? 7'h0 : _GEN_696; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_698 = 10'h2a4 == tempCurrentBuf ? 7'h0 : _GEN_697; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_699 = 10'h2a5 == tempCurrentBuf ? 7'h0 : _GEN_698; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_700 = 10'h2a6 == tempCurrentBuf ? 7'h0 : _GEN_699; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_701 = 10'h2a7 == tempCurrentBuf ? 7'h0 : _GEN_700; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_702 = 10'h2a8 == tempCurrentBuf ? 7'h0 : _GEN_701; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_703 = 10'h2a9 == tempCurrentBuf ? 7'h0 : _GEN_702; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_704 = 10'h2aa == tempCurrentBuf ? 7'h0 : _GEN_703; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_705 = 10'h2ab == tempCurrentBuf ? 7'h0 : _GEN_704; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_706 = 10'h2ac == tempCurrentBuf ? 7'h0 : _GEN_705; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_707 = 10'h2ad == tempCurrentBuf ? 7'h0 : _GEN_706; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_708 = 10'h2ae == tempCurrentBuf ? 7'h0 : _GEN_707; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_709 = 10'h2af == tempCurrentBuf ? 7'h0 : _GEN_708; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_710 = 10'h2b0 == tempCurrentBuf ? 7'h0 : _GEN_709; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_711 = 10'h2b1 == tempCurrentBuf ? 7'h0 : _GEN_710; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_712 = 10'h2b2 == tempCurrentBuf ? 7'h0 : _GEN_711; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_713 = 10'h2b3 == tempCurrentBuf ? 7'h0 : _GEN_712; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_714 = 10'h2b4 == tempCurrentBuf ? 7'h0 : _GEN_713; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_715 = 10'h2b5 == tempCurrentBuf ? 7'h0 : _GEN_714; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_716 = 10'h2b6 == tempCurrentBuf ? 7'h0 : _GEN_715; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_717 = 10'h2b7 == tempCurrentBuf ? 7'h0 : _GEN_716; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_718 = 10'h2b8 == tempCurrentBuf ? 7'h0 : _GEN_717; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_719 = 10'h2b9 == tempCurrentBuf ? 7'h0 : _GEN_718; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_720 = 10'h2ba == tempCurrentBuf ? 7'h0 : _GEN_719; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_721 = 10'h2bb == tempCurrentBuf ? 7'h0 : _GEN_720; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_722 = 10'h2bc == tempCurrentBuf ? 7'h0 : _GEN_721; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_723 = 10'h2bd == tempCurrentBuf ? 7'h0 : _GEN_722; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_724 = 10'h2be == tempCurrentBuf ? 7'h0 : _GEN_723; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_725 = 10'h2bf == tempCurrentBuf ? 7'h0 : _GEN_724; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_726 = 10'h2c0 == tempCurrentBuf ? 7'h0 : _GEN_725; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_727 = 10'h2c1 == tempCurrentBuf ? 7'h0 : _GEN_726; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_728 = 10'h2c2 == tempCurrentBuf ? 7'h0 : _GEN_727; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_729 = 10'h2c3 == tempCurrentBuf ? 7'h0 : _GEN_728; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_730 = 10'h2c4 == tempCurrentBuf ? 7'h0 : _GEN_729; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_731 = 10'h2c5 == tempCurrentBuf ? 7'h0 : _GEN_730; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_732 = 10'h2c6 == tempCurrentBuf ? 7'h0 : _GEN_731; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_733 = 10'h2c7 == tempCurrentBuf ? 7'h0 : _GEN_732; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_734 = 10'h2c8 == tempCurrentBuf ? 7'h0 : _GEN_733; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_735 = 10'h2c9 == tempCurrentBuf ? 7'h0 : _GEN_734; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_736 = 10'h2ca == tempCurrentBuf ? 7'h0 : _GEN_735; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_737 = 10'h2cb == tempCurrentBuf ? 7'h0 : _GEN_736; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_738 = 10'h2cc == tempCurrentBuf ? 7'h0 : _GEN_737; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_739 = 10'h2cd == tempCurrentBuf ? 7'h0 : _GEN_738; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_740 = 10'h2ce == tempCurrentBuf ? 7'h0 : _GEN_739; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_741 = 10'h2cf == tempCurrentBuf ? 7'h0 : _GEN_740; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_742 = 10'h2d0 == tempCurrentBuf ? 7'h0 : _GEN_741; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_743 = 10'h2d1 == tempCurrentBuf ? 7'h0 : _GEN_742; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_744 = 10'h2d2 == tempCurrentBuf ? 7'h0 : _GEN_743; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_745 = 10'h2d3 == tempCurrentBuf ? 7'h0 : _GEN_744; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_746 = 10'h2d4 == tempCurrentBuf ? 7'h0 : _GEN_745; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_747 = 10'h2d5 == tempCurrentBuf ? 7'h0 : _GEN_746; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_748 = 10'h2d6 == tempCurrentBuf ? 7'h0 : _GEN_747; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_749 = 10'h2d7 == tempCurrentBuf ? 7'h0 : _GEN_748; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_750 = 10'h2d8 == tempCurrentBuf ? 7'h0 : _GEN_749; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_751 = 10'h2d9 == tempCurrentBuf ? 7'h0 : _GEN_750; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_752 = 10'h2da == tempCurrentBuf ? 7'h0 : _GEN_751; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_753 = 10'h2db == tempCurrentBuf ? 7'h0 : _GEN_752; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_754 = 10'h2dc == tempCurrentBuf ? 7'h0 : _GEN_753; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_755 = 10'h2dd == tempCurrentBuf ? 7'h0 : _GEN_754; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_756 = 10'h2de == tempCurrentBuf ? 7'h0 : _GEN_755; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_757 = 10'h2df == tempCurrentBuf ? 7'h0 : _GEN_756; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_758 = 10'h2e0 == tempCurrentBuf ? 7'h0 : _GEN_757; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_759 = 10'h2e1 == tempCurrentBuf ? 7'h0 : _GEN_758; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_760 = 10'h2e2 == tempCurrentBuf ? 7'h0 : _GEN_759; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_761 = 10'h2e3 == tempCurrentBuf ? 7'h0 : _GEN_760; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_762 = 10'h2e4 == tempCurrentBuf ? 7'h0 : _GEN_761; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_763 = 10'h2e5 == tempCurrentBuf ? 7'h0 : _GEN_762; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_764 = 10'h2e6 == tempCurrentBuf ? 7'h0 : _GEN_763; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_765 = 10'h2e7 == tempCurrentBuf ? 7'h0 : _GEN_764; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_766 = 10'h2e8 == tempCurrentBuf ? 7'h0 : _GEN_765; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_767 = 10'h2e9 == tempCurrentBuf ? 7'h0 : _GEN_766; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_768 = 10'h2ea == tempCurrentBuf ? 7'h0 : _GEN_767; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_769 = 10'h2eb == tempCurrentBuf ? 7'h0 : _GEN_768; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_770 = 10'h2ec == tempCurrentBuf ? 7'h0 : _GEN_769; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_771 = 10'h2ed == tempCurrentBuf ? 7'h0 : _GEN_770; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_772 = 10'h2ee == tempCurrentBuf ? 7'h0 : _GEN_771; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_773 = 10'h2ef == tempCurrentBuf ? 7'h0 : _GEN_772; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_774 = 10'h2f0 == tempCurrentBuf ? 7'h0 : _GEN_773; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_775 = 10'h2f1 == tempCurrentBuf ? 7'h0 : _GEN_774; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_776 = 10'h2f2 == tempCurrentBuf ? 7'h0 : _GEN_775; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_777 = 10'h2f3 == tempCurrentBuf ? 7'h0 : _GEN_776; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_778 = 10'h2f4 == tempCurrentBuf ? 7'h0 : _GEN_777; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_779 = 10'h2f5 == tempCurrentBuf ? 7'h0 : _GEN_778; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_780 = 10'h2f6 == tempCurrentBuf ? 7'h0 : _GEN_779; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_781 = 10'h2f7 == tempCurrentBuf ? 7'h0 : _GEN_780; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_782 = 10'h2f8 == tempCurrentBuf ? 7'h0 : _GEN_781; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_783 = 10'h2f9 == tempCurrentBuf ? 7'h0 : _GEN_782; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_784 = 10'h2fa == tempCurrentBuf ? 7'h0 : _GEN_783; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_785 = 10'h2fb == tempCurrentBuf ? 7'h0 : _GEN_784; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_786 = 10'h2fc == tempCurrentBuf ? 7'h0 : _GEN_785; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_787 = 10'h2fd == tempCurrentBuf ? 7'h0 : _GEN_786; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_788 = 10'h2fe == tempCurrentBuf ? 7'h0 : _GEN_787; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_789 = 10'h2ff == tempCurrentBuf ? 7'h0 : _GEN_788; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_790 = 10'h300 == tempCurrentBuf ? 7'h0 : _GEN_789; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_791 = 10'h301 == tempCurrentBuf ? 7'h0 : _GEN_790; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_792 = 10'h302 == tempCurrentBuf ? 7'h0 : _GEN_791; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_793 = 10'h303 == tempCurrentBuf ? 7'h0 : _GEN_792; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_794 = 10'h304 == tempCurrentBuf ? 7'h0 : _GEN_793; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_795 = 10'h305 == tempCurrentBuf ? 7'h0 : _GEN_794; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_796 = 10'h306 == tempCurrentBuf ? 7'h0 : _GEN_795; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_797 = 10'h307 == tempCurrentBuf ? 7'h0 : _GEN_796; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_798 = 10'h308 == tempCurrentBuf ? 7'h0 : _GEN_797; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_799 = 10'h309 == tempCurrentBuf ? 7'h0 : _GEN_798; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_800 = 10'h30a == tempCurrentBuf ? 7'h0 : _GEN_799; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_801 = 10'h30b == tempCurrentBuf ? 7'h0 : _GEN_800; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_802 = 10'h30c == tempCurrentBuf ? 7'h0 : _GEN_801; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_803 = 10'h30d == tempCurrentBuf ? 7'h0 : _GEN_802; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_804 = 10'h30e == tempCurrentBuf ? 7'h0 : _GEN_803; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_805 = 10'h30f == tempCurrentBuf ? 7'h0 : _GEN_804; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_806 = 10'h310 == tempCurrentBuf ? 7'h0 : _GEN_805; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_807 = 10'h311 == tempCurrentBuf ? 7'h0 : _GEN_806; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_808 = 10'h312 == tempCurrentBuf ? 7'h0 : _GEN_807; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_809 = 10'h313 == tempCurrentBuf ? 7'h0 : _GEN_808; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_810 = 10'h314 == tempCurrentBuf ? 7'h0 : _GEN_809; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_811 = 10'h315 == tempCurrentBuf ? 7'h0 : _GEN_810; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_812 = 10'h316 == tempCurrentBuf ? 7'h0 : _GEN_811; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_813 = 10'h317 == tempCurrentBuf ? 7'h0 : _GEN_812; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_814 = 10'h318 == tempCurrentBuf ? 7'h0 : _GEN_813; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_815 = 10'h319 == tempCurrentBuf ? 7'h0 : _GEN_814; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_816 = 10'h31a == tempCurrentBuf ? 7'h0 : _GEN_815; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_817 = 10'h31b == tempCurrentBuf ? 7'h0 : _GEN_816; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_818 = 10'h31c == tempCurrentBuf ? 7'h0 : _GEN_817; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_819 = 10'h31d == tempCurrentBuf ? 7'h0 : _GEN_818; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_820 = 10'h31e == tempCurrentBuf ? 7'h0 : _GEN_819; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_821 = 10'h31f == tempCurrentBuf ? 7'h0 : _GEN_820; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_822 = 10'h320 == tempCurrentBuf ? 7'h0 : _GEN_821; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_823 = 10'h321 == tempCurrentBuf ? 7'h0 : _GEN_822; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_824 = 10'h322 == tempCurrentBuf ? 7'h0 : _GEN_823; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_825 = 10'h323 == tempCurrentBuf ? 7'h0 : _GEN_824; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_826 = 10'h324 == tempCurrentBuf ? 7'h0 : _GEN_825; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_827 = 10'h325 == tempCurrentBuf ? 7'h0 : _GEN_826; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_828 = 10'h326 == tempCurrentBuf ? 7'h0 : _GEN_827; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_829 = 10'h327 == tempCurrentBuf ? 7'h0 : _GEN_828; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_830 = 10'h328 == tempCurrentBuf ? 7'h0 : _GEN_829; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_831 = 10'h329 == tempCurrentBuf ? 7'h0 : _GEN_830; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_832 = 10'h32a == tempCurrentBuf ? 7'h0 : _GEN_831; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_833 = 10'h32b == tempCurrentBuf ? 7'h0 : _GEN_832; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_834 = 10'h32c == tempCurrentBuf ? 7'h0 : _GEN_833; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_835 = 10'h32d == tempCurrentBuf ? 7'h0 : _GEN_834; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_836 = 10'h32e == tempCurrentBuf ? 7'h0 : _GEN_835; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_837 = 10'h32f == tempCurrentBuf ? 7'h0 : _GEN_836; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_838 = 10'h330 == tempCurrentBuf ? 7'h0 : _GEN_837; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_839 = 10'h331 == tempCurrentBuf ? 7'h0 : _GEN_838; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_840 = 10'h332 == tempCurrentBuf ? 7'h0 : _GEN_839; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_841 = 10'h333 == tempCurrentBuf ? 7'h0 : _GEN_840; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_842 = 10'h334 == tempCurrentBuf ? 7'h0 : _GEN_841; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_843 = 10'h335 == tempCurrentBuf ? 7'h0 : _GEN_842; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_844 = 10'h336 == tempCurrentBuf ? 7'h0 : _GEN_843; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_845 = 10'h337 == tempCurrentBuf ? 7'h0 : _GEN_844; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_846 = 10'h338 == tempCurrentBuf ? 7'h0 : _GEN_845; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_847 = 10'h339 == tempCurrentBuf ? 7'h0 : _GEN_846; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_848 = 10'h33a == tempCurrentBuf ? 7'h0 : _GEN_847; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_849 = 10'h33b == tempCurrentBuf ? 7'h0 : _GEN_848; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_850 = 10'h33c == tempCurrentBuf ? 7'h0 : _GEN_849; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_851 = 10'h33d == tempCurrentBuf ? 7'h0 : _GEN_850; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_852 = 10'h33e == tempCurrentBuf ? 7'h0 : _GEN_851; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_853 = 10'h33f == tempCurrentBuf ? 7'h0 : _GEN_852; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_854 = 10'h340 == tempCurrentBuf ? 7'h0 : _GEN_853; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_855 = 10'h341 == tempCurrentBuf ? 7'h0 : _GEN_854; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_856 = 10'h342 == tempCurrentBuf ? 7'h0 : _GEN_855; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_857 = 10'h343 == tempCurrentBuf ? 7'h0 : _GEN_856; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_858 = 10'h344 == tempCurrentBuf ? 7'h0 : _GEN_857; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_859 = 10'h345 == tempCurrentBuf ? 7'h0 : _GEN_858; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_860 = 10'h346 == tempCurrentBuf ? 7'h0 : _GEN_859; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_861 = 10'h347 == tempCurrentBuf ? 7'h0 : _GEN_860; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_862 = 10'h348 == tempCurrentBuf ? 7'h0 : _GEN_861; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_863 = 10'h349 == tempCurrentBuf ? 7'h0 : _GEN_862; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_864 = 10'h34a == tempCurrentBuf ? 7'h0 : _GEN_863; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_865 = 10'h34b == tempCurrentBuf ? 7'h0 : _GEN_864; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_866 = 10'h34c == tempCurrentBuf ? 7'h0 : _GEN_865; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_867 = 10'h34d == tempCurrentBuf ? 7'h0 : _GEN_866; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_868 = 10'h34e == tempCurrentBuf ? 7'h0 : _GEN_867; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_869 = 10'h34f == tempCurrentBuf ? 7'h0 : _GEN_868; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_870 = 10'h350 == tempCurrentBuf ? 7'h0 : _GEN_869; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_871 = 10'h351 == tempCurrentBuf ? 7'h0 : _GEN_870; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_872 = 10'h352 == tempCurrentBuf ? 7'h0 : _GEN_871; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_873 = 10'h353 == tempCurrentBuf ? 7'h0 : _GEN_872; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_874 = 10'h354 == tempCurrentBuf ? 7'h0 : _GEN_873; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_875 = 10'h355 == tempCurrentBuf ? 7'h0 : _GEN_874; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_876 = 10'h356 == tempCurrentBuf ? 7'h0 : _GEN_875; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_877 = 10'h357 == tempCurrentBuf ? 7'h0 : _GEN_876; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_878 = 10'h358 == tempCurrentBuf ? 7'h0 : _GEN_877; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_879 = 10'h359 == tempCurrentBuf ? 7'h0 : _GEN_878; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_880 = 10'h35a == tempCurrentBuf ? 7'h0 : _GEN_879; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_881 = 10'h35b == tempCurrentBuf ? 7'h0 : _GEN_880; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_882 = 10'h35c == tempCurrentBuf ? 7'h0 : _GEN_881; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_883 = 10'h35d == tempCurrentBuf ? 7'h0 : _GEN_882; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_884 = 10'h35e == tempCurrentBuf ? 7'h0 : _GEN_883; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_885 = 10'h35f == tempCurrentBuf ? 7'h0 : _GEN_884; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_886 = 10'h360 == tempCurrentBuf ? 7'h0 : _GEN_885; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_887 = 10'h361 == tempCurrentBuf ? 7'h0 : _GEN_886; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_888 = 10'h362 == tempCurrentBuf ? 7'h0 : _GEN_887; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_889 = 10'h363 == tempCurrentBuf ? 7'h0 : _GEN_888; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_890 = 10'h364 == tempCurrentBuf ? 7'h0 : _GEN_889; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_891 = 10'h365 == tempCurrentBuf ? 7'h0 : _GEN_890; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_892 = 10'h366 == tempCurrentBuf ? 7'h0 : _GEN_891; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_893 = 10'h367 == tempCurrentBuf ? 7'h0 : _GEN_892; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_894 = 10'h368 == tempCurrentBuf ? 7'h0 : _GEN_893; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_895 = 10'h369 == tempCurrentBuf ? 7'h0 : _GEN_894; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_896 = 10'h36a == tempCurrentBuf ? 7'h0 : _GEN_895; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_897 = 10'h36b == tempCurrentBuf ? 7'h0 : _GEN_896; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_898 = 10'h36c == tempCurrentBuf ? 7'h0 : _GEN_897; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_899 = 10'h36d == tempCurrentBuf ? 7'h0 : _GEN_898; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_900 = 10'h36e == tempCurrentBuf ? 7'h0 : _GEN_899; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_901 = 10'h36f == tempCurrentBuf ? 7'h0 : _GEN_900; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_902 = 10'h370 == tempCurrentBuf ? 7'h0 : _GEN_901; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_903 = 10'h371 == tempCurrentBuf ? 7'h0 : _GEN_902; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_904 = 10'h372 == tempCurrentBuf ? 7'h0 : _GEN_903; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_905 = 10'h373 == tempCurrentBuf ? 7'h0 : _GEN_904; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_906 = 10'h374 == tempCurrentBuf ? 7'h0 : _GEN_905; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_907 = 10'h375 == tempCurrentBuf ? 7'h0 : _GEN_906; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_908 = 10'h376 == tempCurrentBuf ? 7'h0 : _GEN_907; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_909 = 10'h377 == tempCurrentBuf ? 7'h0 : _GEN_908; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_910 = 10'h378 == tempCurrentBuf ? 7'h0 : _GEN_909; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_911 = 10'h379 == tempCurrentBuf ? 7'h0 : _GEN_910; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_912 = 10'h37a == tempCurrentBuf ? 7'h0 : _GEN_911; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_913 = 10'h37b == tempCurrentBuf ? 7'h0 : _GEN_912; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_914 = 10'h37c == tempCurrentBuf ? 7'h0 : _GEN_913; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_915 = 10'h37d == tempCurrentBuf ? 7'h0 : _GEN_914; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_916 = 10'h37e == tempCurrentBuf ? 7'h0 : _GEN_915; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_917 = 10'h37f == tempCurrentBuf ? 7'h0 : _GEN_916; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_918 = 10'h380 == tempCurrentBuf ? 7'h0 : _GEN_917; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_919 = 10'h381 == tempCurrentBuf ? 7'h0 : _GEN_918; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_920 = 10'h382 == tempCurrentBuf ? 7'h0 : _GEN_919; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_921 = 10'h383 == tempCurrentBuf ? 7'h0 : _GEN_920; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_922 = 10'h384 == tempCurrentBuf ? 7'h0 : _GEN_921; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_923 = 10'h385 == tempCurrentBuf ? 7'h0 : _GEN_922; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_924 = 10'h386 == tempCurrentBuf ? 7'h0 : _GEN_923; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_925 = 10'h387 == tempCurrentBuf ? 7'h0 : _GEN_924; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_926 = 10'h388 == tempCurrentBuf ? 7'h0 : _GEN_925; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_927 = 10'h389 == tempCurrentBuf ? 7'h0 : _GEN_926; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_928 = 10'h38a == tempCurrentBuf ? 7'h0 : _GEN_927; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_929 = 10'h38b == tempCurrentBuf ? 7'h0 : _GEN_928; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_930 = 10'h38c == tempCurrentBuf ? 7'h0 : _GEN_929; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_931 = 10'h38d == tempCurrentBuf ? 7'h0 : _GEN_930; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_932 = 10'h38e == tempCurrentBuf ? 7'h0 : _GEN_931; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_933 = 10'h38f == tempCurrentBuf ? 7'h0 : _GEN_932; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_934 = 10'h390 == tempCurrentBuf ? 7'h0 : _GEN_933; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_935 = 10'h391 == tempCurrentBuf ? 7'h0 : _GEN_934; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_936 = 10'h392 == tempCurrentBuf ? 7'h0 : _GEN_935; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_937 = 10'h393 == tempCurrentBuf ? 7'h0 : _GEN_936; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_938 = 10'h394 == tempCurrentBuf ? 7'h0 : _GEN_937; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_939 = 10'h395 == tempCurrentBuf ? 7'h0 : _GEN_938; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_940 = 10'h396 == tempCurrentBuf ? 7'h0 : _GEN_939; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_941 = 10'h397 == tempCurrentBuf ? 7'h0 : _GEN_940; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_942 = 10'h398 == tempCurrentBuf ? 7'h0 : _GEN_941; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_943 = 10'h399 == tempCurrentBuf ? 7'h0 : _GEN_942; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_944 = 10'h39a == tempCurrentBuf ? 7'h0 : _GEN_943; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_945 = 10'h39b == tempCurrentBuf ? 7'h0 : _GEN_944; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_946 = 10'h39c == tempCurrentBuf ? 7'h0 : _GEN_945; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_947 = 10'h39d == tempCurrentBuf ? 7'h0 : _GEN_946; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_948 = 10'h39e == tempCurrentBuf ? 7'h0 : _GEN_947; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_949 = 10'h39f == tempCurrentBuf ? 7'h0 : _GEN_948; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_950 = 10'h3a0 == tempCurrentBuf ? 7'h0 : _GEN_949; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_951 = 10'h3a1 == tempCurrentBuf ? 7'h0 : _GEN_950; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_952 = 10'h3a2 == tempCurrentBuf ? 7'h0 : _GEN_951; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_953 = 10'h3a3 == tempCurrentBuf ? 7'h0 : _GEN_952; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_954 = 10'h3a4 == tempCurrentBuf ? 7'h0 : _GEN_953; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_955 = 10'h3a5 == tempCurrentBuf ? 7'h0 : _GEN_954; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_956 = 10'h3a6 == tempCurrentBuf ? 7'h0 : _GEN_955; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_957 = 10'h3a7 == tempCurrentBuf ? 7'h0 : _GEN_956; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_958 = 10'h3a8 == tempCurrentBuf ? 7'h0 : _GEN_957; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_959 = 10'h3a9 == tempCurrentBuf ? 7'h0 : _GEN_958; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_960 = 10'h3aa == tempCurrentBuf ? 7'h0 : _GEN_959; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_961 = 10'h3ab == tempCurrentBuf ? 7'h0 : _GEN_960; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_962 = 10'h3ac == tempCurrentBuf ? 7'h0 : _GEN_961; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_963 = 10'h3ad == tempCurrentBuf ? 7'h0 : _GEN_962; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_964 = 10'h3ae == tempCurrentBuf ? 7'h0 : _GEN_963; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_965 = 10'h3af == tempCurrentBuf ? 7'h0 : _GEN_964; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_966 = 10'h3b0 == tempCurrentBuf ? 7'h0 : _GEN_965; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_967 = 10'h3b1 == tempCurrentBuf ? 7'h0 : _GEN_966; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_968 = 10'h3b2 == tempCurrentBuf ? 7'h0 : _GEN_967; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_969 = 10'h3b3 == tempCurrentBuf ? 7'h0 : _GEN_968; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_970 = 10'h3b4 == tempCurrentBuf ? 7'h0 : _GEN_969; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_971 = 10'h3b5 == tempCurrentBuf ? 7'h0 : _GEN_970; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_972 = 10'h3b6 == tempCurrentBuf ? 7'h0 : _GEN_971; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_973 = 10'h3b7 == tempCurrentBuf ? 7'h0 : _GEN_972; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_974 = 10'h3b8 == tempCurrentBuf ? 7'h0 : _GEN_973; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_975 = 10'h3b9 == tempCurrentBuf ? 7'h0 : _GEN_974; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_976 = 10'h3ba == tempCurrentBuf ? 7'h0 : _GEN_975; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_977 = 10'h3bb == tempCurrentBuf ? 7'h0 : _GEN_976; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_978 = 10'h3bc == tempCurrentBuf ? 7'h0 : _GEN_977; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_979 = 10'h3bd == tempCurrentBuf ? 7'h0 : _GEN_978; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_980 = 10'h3be == tempCurrentBuf ? 7'h0 : _GEN_979; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_981 = 10'h3bf == tempCurrentBuf ? 7'h0 : _GEN_980; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_982 = 10'h3c0 == tempCurrentBuf ? 7'h0 : _GEN_981; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_983 = 10'h3c1 == tempCurrentBuf ? 7'h0 : _GEN_982; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_984 = 10'h3c2 == tempCurrentBuf ? 7'h0 : _GEN_983; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_985 = 10'h3c3 == tempCurrentBuf ? 7'h0 : _GEN_984; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_986 = 10'h3c4 == tempCurrentBuf ? 7'h0 : _GEN_985; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_987 = 10'h3c5 == tempCurrentBuf ? 7'h0 : _GEN_986; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_988 = 10'h3c6 == tempCurrentBuf ? 7'h0 : _GEN_987; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_989 = 10'h3c7 == tempCurrentBuf ? 7'h0 : _GEN_988; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_990 = 10'h3c8 == tempCurrentBuf ? 7'h0 : _GEN_989; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_991 = 10'h3c9 == tempCurrentBuf ? 7'h0 : _GEN_990; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_992 = 10'h3ca == tempCurrentBuf ? 7'h0 : _GEN_991; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_993 = 10'h3cb == tempCurrentBuf ? 7'h0 : _GEN_992; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_994 = 10'h3cc == tempCurrentBuf ? 7'h0 : _GEN_993; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_995 = 10'h3cd == tempCurrentBuf ? 7'h0 : _GEN_994; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_996 = 10'h3ce == tempCurrentBuf ? 7'h0 : _GEN_995; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_997 = 10'h3cf == tempCurrentBuf ? 7'h0 : _GEN_996; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_998 = 10'h3d0 == tempCurrentBuf ? 7'h0 : _GEN_997; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_999 = 10'h3d1 == tempCurrentBuf ? 7'h0 : _GEN_998; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1000 = 10'h3d2 == tempCurrentBuf ? 7'h0 : _GEN_999; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1001 = 10'h3d3 == tempCurrentBuf ? 7'h0 : _GEN_1000; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1002 = 10'h3d4 == tempCurrentBuf ? 7'h0 : _GEN_1001; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1003 = 10'h3d5 == tempCurrentBuf ? 7'h0 : _GEN_1002; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1004 = 10'h3d6 == tempCurrentBuf ? 7'h0 : _GEN_1003; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1005 = 10'h3d7 == tempCurrentBuf ? 7'h0 : _GEN_1004; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1006 = 10'h3d8 == tempCurrentBuf ? 7'h0 : _GEN_1005; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1007 = 10'h3d9 == tempCurrentBuf ? 7'h0 : _GEN_1006; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1008 = 10'h3da == tempCurrentBuf ? 7'h0 : _GEN_1007; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1009 = 10'h3db == tempCurrentBuf ? 7'h0 : _GEN_1008; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1010 = 10'h3dc == tempCurrentBuf ? 7'h0 : _GEN_1009; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1011 = 10'h3dd == tempCurrentBuf ? 7'h0 : _GEN_1010; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1012 = 10'h3de == tempCurrentBuf ? 7'h0 : _GEN_1011; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1013 = 10'h3df == tempCurrentBuf ? 7'h0 : _GEN_1012; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1014 = 10'h3e0 == tempCurrentBuf ? 7'h0 : _GEN_1013; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1015 = 10'h3e1 == tempCurrentBuf ? 7'h0 : _GEN_1014; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1016 = 10'h3e2 == tempCurrentBuf ? 7'h0 : _GEN_1015; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1017 = 10'h3e3 == tempCurrentBuf ? 7'h0 : _GEN_1016; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1018 = 10'h3e4 == tempCurrentBuf ? 7'h0 : _GEN_1017; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1019 = 10'h3e5 == tempCurrentBuf ? 7'h0 : _GEN_1018; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1020 = 10'h3e6 == tempCurrentBuf ? 7'h0 : _GEN_1019; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1021 = 10'h3e7 == tempCurrentBuf ? 7'h0 : _GEN_1020; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1022 = 10'h3e8 == tempCurrentBuf ? 7'h0 : _GEN_1021; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1023 = 10'h3e9 == tempCurrentBuf ? 7'h0 : _GEN_1022; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1024 = 10'h3ea == tempCurrentBuf ? 7'h0 : _GEN_1023; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1025 = 10'h3eb == tempCurrentBuf ? 7'h0 : _GEN_1024; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1026 = 10'h3ec == tempCurrentBuf ? 7'h0 : _GEN_1025; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1027 = 10'h3ed == tempCurrentBuf ? 7'h0 : _GEN_1026; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1028 = 10'h3ee == tempCurrentBuf ? 7'h0 : _GEN_1027; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1029 = 10'h3ef == tempCurrentBuf ? 7'h0 : _GEN_1028; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1030 = 10'h3f0 == tempCurrentBuf ? 7'h0 : _GEN_1029; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1031 = 10'h3f1 == tempCurrentBuf ? 7'h0 : _GEN_1030; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1032 = 10'h3f2 == tempCurrentBuf ? 7'h0 : _GEN_1031; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1033 = 10'h3f3 == tempCurrentBuf ? 7'h0 : _GEN_1032; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1034 = 10'h3f4 == tempCurrentBuf ? 7'h0 : _GEN_1033; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1035 = 10'h3f5 == tempCurrentBuf ? 7'h0 : _GEN_1034; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1036 = 10'h3f6 == tempCurrentBuf ? 7'h0 : _GEN_1035; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1037 = 10'h3f7 == tempCurrentBuf ? 7'h0 : _GEN_1036; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1038 = 10'h3f8 == tempCurrentBuf ? 7'h0 : _GEN_1037; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1039 = 10'h3f9 == tempCurrentBuf ? 7'h0 : _GEN_1038; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1040 = 10'h3fa == tempCurrentBuf ? 7'h0 : _GEN_1039; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1041 = 10'h3fb == tempCurrentBuf ? 7'h0 : _GEN_1040; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1042 = 10'h3fc == tempCurrentBuf ? 7'h0 : _GEN_1041; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1043 = 10'h3fd == tempCurrentBuf ? 7'h0 : _GEN_1042; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1044 = 10'h3fe == tempCurrentBuf ? 7'h0 : _GEN_1043; // @[lut_mem_online2.scala 148:{24,24}]
  wire [6:0] _GEN_1045 = 10'h3ff == tempCurrentBuf ? 7'h0 : _GEN_1044; // @[lut_mem_online2.scala 148:{24,24}]
  wire [3:0] _outResult_T_1 = 4'h6 - outputCounter; // @[lut_mem_online2.scala 165:60]
  wire [6:0] _outResult_T_2 = outputBuffer >> _outResult_T_1; // @[lut_mem_online2.scala 165:36]
  wire [3:0] _outputCounter_T_1 = outputCounter + 4'h1; // @[lut_mem_online2.scala 167:42]
  wire  _GEN_1047 = isOutputValid & outputCounter != 4'h7 & _outResult_T_2[0]; // @[lut_mem_online2.scala 163:78 165:21 172:23]
  assign io_outResult = outResult; // @[lut_mem_online2.scala 209:16]
  always @(posedge clock) begin
    buffer_0 <= io_start & _GEN_11; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_1 <= io_start & _GEN_12; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_2 <= io_start & _GEN_13; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_3 <= io_start & _GEN_14; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_4 <= io_start & _GEN_15; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_5 <= io_start & _GEN_16; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_6 <= io_start & _GEN_17; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_7 <= io_start & _GEN_18; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_8 <= io_start & _GEN_19; // @[lut_mem_online2.scala 198:17 98:29]
    buffer_9 <= io_start & _GEN_20; // @[lut_mem_online2.scala 198:17 98:29]
    if (reset) begin // @[lut_mem_online2.scala 77:29]
      outputBuffer <= 7'h0; // @[lut_mem_online2.scala 77:29]
    end else if (io_start) begin // @[lut_mem_online2.scala 98:29]
      if (isPassedDelta) begin // @[lut_mem_online2.scala 143:40]
        if (10'h3ff == tempCurrentBuf) begin // @[lut_mem_online2.scala 148:24]
          outputBuffer <= 7'h0; // @[lut_mem_online2.scala 148:24]
        end else begin
          outputBuffer <= _GEN_1044;
        end
      end
    end
    if (reset) begin // @[lut_mem_online2.scala 79:24]
      counter <= 4'h0; // @[lut_mem_online2.scala 79:24]
    end else if (io_start) begin // @[lut_mem_online2.scala 98:29]
      if (counter != 4'ha) begin // @[lut_mem_online2.scala 121:38]
        counter <= _counter_T_1; // @[lut_mem_online2.scala 137:19]
      end
    end else begin
      counter <= 4'h0; // @[lut_mem_online2.scala 194:13]
    end
    if (reset) begin // @[lut_mem_online2.scala 80:30]
      outputCounter <= 4'h0; // @[lut_mem_online2.scala 80:30]
    end else if (io_start) begin // @[lut_mem_online2.scala 98:29]
      if (isOutputValid & outputCounter != 4'h7) begin // @[lut_mem_online2.scala 163:78]
        outputCounter <= _outputCounter_T_1; // @[lut_mem_online2.scala 167:25]
      end
    end else begin
      outputCounter <= 4'h0; // @[lut_mem_online2.scala 195:19]
    end
    if (reset) begin // @[lut_mem_online2.scala 82:30]
      isPassedDelta <= 1'h0; // @[lut_mem_online2.scala 82:30]
    end else if (io_start) begin // @[lut_mem_online2.scala 98:29]
      isPassedDelta <= _GEN_0;
    end
    isOutputValid <= isPassedDelta; // @[lut_mem_online2.scala 83:30]
    if (reset) begin // @[lut_mem_online2.scala 86:26]
      outResult <= 1'h0; // @[lut_mem_online2.scala 86:26]
    end else if (io_start) begin // @[lut_mem_online2.scala 98:29]
      outResult <= _GEN_1047;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_3 & ~reset) begin
          $fwrite(32'h80000002,"buffer(%d) = %d\n",counter,io_inputBit); // @[lut_mem_online2.scala 127:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & isPassedDelta & _T_5) begin
          $fwrite(32'h80000002,"lut(%d) = %d\n",tempCurrentBuf,_GEN_1045); // @[lut_mem_online2.scala 152:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
