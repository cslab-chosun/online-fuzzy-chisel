module LutMembershipFunctionOnline_3(
  input   clock,
  input   reset,
  input   io_start,
  input   io_inputBit,
  output  io_outResult
);
  reg [7:0] i; // @[lut_mem_online.scala 205:18]
  reg  buffer_0; // @[lut_mem_online.scala 209:19]
  reg  buffer_1; // @[lut_mem_online.scala 209:19]
  reg  buffer_2; // @[lut_mem_online.scala 209:19]
  reg  buffer_3; // @[lut_mem_online.scala 209:19]
  reg  buffer_4; // @[lut_mem_online.scala 209:19]
  reg  buffer_5; // @[lut_mem_online.scala 209:19]
  reg  buffer_6; // @[lut_mem_online.scala 209:19]
  reg [3:0] counter; // @[lut_mem_online.scala 211:24]
  reg  outResult; // @[lut_mem_online.scala 214:26]
  wire  _T_2 = counter < 4'h8; // @[lut_mem_online.scala 231:22]
  wire  _GEN_0 = io_inputBit ? 1'h0 : buffer_0; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_1 = i == 8'h0 ? _GEN_0 : buffer_0; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_2 = io_inputBit ? 1'h0 : _GEN_1; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_3 = i == 8'h1 ? _GEN_2 : _GEN_1; // @[lut_mem_online.scala 234:34]
  wire  _GEN_4 = io_inputBit ? 1'h0 : _GEN_3; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_5 = i == 8'h3 ? _GEN_4 : _GEN_3; // @[lut_mem_online.scala 234:34]
  wire  _T_10 = ~io_inputBit; // @[lut_mem_online.scala 236:32]
  wire  _GEN_6 = ~io_inputBit | _GEN_5; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_7 = i == 8'h7 ? _GEN_6 : _GEN_5; // @[lut_mem_online.scala 234:34]
  wire  _GEN_8 = ~io_inputBit | _GEN_7; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_9 = i == 8'h10 ? _GEN_8 : _GEN_7; // @[lut_mem_online.scala 234:34]
  wire  _GEN_10 = ~io_inputBit | _GEN_9; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_11 = i == 8'h22 ? _GEN_10 : _GEN_9; // @[lut_mem_online.scala 234:34]
  wire  _GEN_12 = io_inputBit ? 1'h0 : _GEN_11; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_13 = i == 8'h22 ? _GEN_12 : _GEN_11; // @[lut_mem_online.scala 234:34]
  wire  _GEN_14 = io_inputBit ? 1'h0 : buffer_1; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_15 = i == 8'h0 ? _GEN_14 : buffer_1; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_16 = io_inputBit ? 1'h0 : _GEN_15; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_17 = i == 8'h1 ? _GEN_16 : _GEN_15; // @[lut_mem_online.scala 234:34]
  wire  _GEN_18 = ~io_inputBit | _GEN_17; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_19 = i == 8'h7 ? _GEN_18 : _GEN_17; // @[lut_mem_online.scala 234:34]
  wire  _GEN_20 = io_inputBit ? 1'h0 : _GEN_19; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_21 = i == 8'h8 ? _GEN_20 : _GEN_19; // @[lut_mem_online.scala 234:34]
  wire  _GEN_22 = io_inputBit ? 1'h0 : _GEN_21; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_23 = i == 8'h11 ? _GEN_22 : _GEN_21; // @[lut_mem_online.scala 234:34]
  wire  _GEN_24 = ~io_inputBit | _GEN_23; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_25 = i == 8'h21 ? _GEN_24 : _GEN_23; // @[lut_mem_online.scala 234:34]
  wire  _GEN_26 = ~io_inputBit ? 1'h0 : _GEN_25; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_27 = i == 8'h22 ? _GEN_26 : _GEN_25; // @[lut_mem_online.scala 234:34]
  wire  _GEN_28 = io_inputBit | _GEN_27; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_29 = i == 8'h22 ? _GEN_28 : _GEN_27; // @[lut_mem_online.scala 234:34]
  wire  _GEN_30 = io_inputBit ? 1'h0 : _GEN_29; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_31 = i == 8'h23 ? _GEN_30 : _GEN_29; // @[lut_mem_online.scala 234:34]
  wire  _GEN_32 = io_inputBit ? 1'h0 : _GEN_31; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_33 = i == 8'h44 ? _GEN_32 : _GEN_31; // @[lut_mem_online.scala 234:34]
  wire  _GEN_34 = ~io_inputBit | _GEN_33; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_35 = i == 8'h47 ? _GEN_34 : _GEN_33; // @[lut_mem_online.scala 234:34]
  wire  _GEN_36 = io_inputBit ? 1'h0 : _GEN_35; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_37 = i == 8'h47 ? _GEN_36 : _GEN_35; // @[lut_mem_online.scala 234:34]
  wire  _GEN_38 = ~io_inputBit | _GEN_37; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_39 = i == 8'h89 ? _GEN_38 : _GEN_37; // @[lut_mem_online.scala 234:34]
  wire  _GEN_40 = io_inputBit ? 1'h0 : _GEN_39; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_41 = i == 8'h89 ? _GEN_40 : _GEN_39; // @[lut_mem_online.scala 234:34]
  wire  _GEN_42 = io_inputBit ? 1'h0 : buffer_2; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_43 = i == 8'h0 ? _GEN_42 : buffer_2; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_44 = io_inputBit ? 1'h0 : _GEN_43; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_45 = i == 8'h1 ? _GEN_44 : _GEN_43; // @[lut_mem_online.scala 234:34]
  wire  _GEN_46 = ~io_inputBit ? 1'h0 : _GEN_45; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_47 = i == 8'h7 ? _GEN_46 : _GEN_45; // @[lut_mem_online.scala 234:34]
  wire  _GEN_48 = io_inputBit ? 1'h0 : _GEN_47; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_49 = i == 8'h8 ? _GEN_48 : _GEN_47; // @[lut_mem_online.scala 234:34]
  wire  _GEN_50 = io_inputBit ? 1'h0 : _GEN_49; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_51 = i == 8'h11 ? _GEN_50 : _GEN_49; // @[lut_mem_online.scala 234:34]
  wire  _GEN_52 = ~io_inputBit ? 1'h0 : _GEN_51; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_53 = i == 8'h21 ? _GEN_52 : _GEN_51; // @[lut_mem_online.scala 234:34]
  wire  _GEN_54 = io_inputBit | _GEN_53; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_55 = i == 8'h44 ? _GEN_54 : _GEN_53; // @[lut_mem_online.scala 234:34]
  wire  _GEN_56 = io_inputBit ? 1'h0 : _GEN_55; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_57 = i == 8'h45 ? _GEN_56 : _GEN_55; // @[lut_mem_online.scala 234:34]
  wire  _GEN_58 = ~io_inputBit | _GEN_57; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_59 = i == 8'h46 ? _GEN_58 : _GEN_57; // @[lut_mem_online.scala 234:34]
  wire  _GEN_60 = ~io_inputBit ? 1'h0 : _GEN_59; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_61 = i == 8'h47 ? _GEN_60 : _GEN_59; // @[lut_mem_online.scala 234:34]
  wire  _GEN_62 = io_inputBit | _GEN_61; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_63 = i == 8'h47 ? _GEN_62 : _GEN_61; // @[lut_mem_online.scala 234:34]
  wire  _GEN_64 = io_inputBit ? 1'h0 : _GEN_63; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_65 = i == 8'h48 ? _GEN_64 : _GEN_63; // @[lut_mem_online.scala 234:34]
  wire  _GEN_66 = ~io_inputBit ? 1'h0 : _GEN_65; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_67 = i == 8'h89 ? _GEN_66 : _GEN_65; // @[lut_mem_online.scala 234:34]
  wire  _GEN_68 = io_inputBit | _GEN_67; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_69 = i == 8'h89 ? _GEN_68 : _GEN_67; // @[lut_mem_online.scala 234:34]
  wire  _GEN_70 = ~io_inputBit | _GEN_69; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_71 = i == 8'h8b ? _GEN_70 : _GEN_69; // @[lut_mem_online.scala 234:34]
  wire  _GEN_72 = io_inputBit ? 1'h0 : _GEN_71; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_73 = i == 8'h8b ? _GEN_72 : _GEN_71; // @[lut_mem_online.scala 234:34]
  wire  _GEN_74 = ~io_inputBit | _GEN_73; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_75 = i == 8'h8e ? _GEN_74 : _GEN_73; // @[lut_mem_online.scala 234:34]
  wire  _GEN_76 = io_inputBit ? 1'h0 : _GEN_75; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_77 = i == 8'h8e ? _GEN_76 : _GEN_75; // @[lut_mem_online.scala 234:34]
  wire  _GEN_78 = ~io_inputBit | _GEN_77; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_79 = i == 8'h91 ? _GEN_78 : _GEN_77; // @[lut_mem_online.scala 234:34]
  wire  _GEN_80 = io_inputBit ? 1'h0 : _GEN_79; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_81 = i == 8'h91 ? _GEN_80 : _GEN_79; // @[lut_mem_online.scala 234:34]
  wire  _GEN_82 = io_inputBit ? 1'h0 : buffer_3; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_83 = i == 8'h0 ? _GEN_82 : buffer_3; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_84 = io_inputBit ? 1'h0 : _GEN_83; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_85 = i == 8'h1 ? _GEN_84 : _GEN_83; // @[lut_mem_online.scala 234:34]
  wire  _GEN_86 = ~io_inputBit ? 1'h0 : _GEN_85; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_87 = i == 8'h7 ? _GEN_86 : _GEN_85; // @[lut_mem_online.scala 234:34]
  wire  _GEN_88 = io_inputBit ? 1'h0 : _GEN_87; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_89 = i == 8'h8 ? _GEN_88 : _GEN_87; // @[lut_mem_online.scala 234:34]
  wire  _GEN_90 = io_inputBit ? 1'h0 : _GEN_89; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_91 = i == 8'h11 ? _GEN_90 : _GEN_89; // @[lut_mem_online.scala 234:34]
  wire  _GEN_92 = ~io_inputBit ? 1'h0 : _GEN_91; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_93 = i == 8'h21 ? _GEN_92 : _GEN_91; // @[lut_mem_online.scala 234:34]
  wire  _GEN_94 = io_inputBit ? 1'h0 : _GEN_93; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_95 = i == 8'h45 ? _GEN_94 : _GEN_93; // @[lut_mem_online.scala 234:34]
  wire  _GEN_96 = io_inputBit | _GEN_95; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_97 = i == 8'h47 ? _GEN_96 : _GEN_95; // @[lut_mem_online.scala 234:34]
  wire  _GEN_98 = ~io_inputBit ? 1'h0 : _GEN_97; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_99 = i == 8'h89 ? _GEN_98 : _GEN_97; // @[lut_mem_online.scala 234:34]
  wire  _GEN_100 = io_inputBit | _GEN_99; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_101 = i == 8'h89 ? _GEN_100 : _GEN_99; // @[lut_mem_online.scala 234:34]
  wire  _GEN_102 = ~io_inputBit | _GEN_101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_103 = i == 8'h8a ? _GEN_102 : _GEN_101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_104 = io_inputBit ? 1'h0 : _GEN_103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_105 = i == 8'h8a ? _GEN_104 : _GEN_103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_106 = ~io_inputBit ? 1'h0 : _GEN_105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_107 = i == 8'h8b ? _GEN_106 : _GEN_105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_108 = io_inputBit | _GEN_107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_109 = i == 8'h8b ? _GEN_108 : _GEN_107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_110 = ~io_inputBit | _GEN_109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_111 = i == 8'h8d ? _GEN_110 : _GEN_109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_112 = io_inputBit ? 1'h0 : _GEN_111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_113 = i == 8'h8d ? _GEN_112 : _GEN_111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_114 = ~io_inputBit ? 1'h0 : _GEN_113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_115 = i == 8'h8e ? _GEN_114 : _GEN_113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_116 = io_inputBit | _GEN_115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_117 = i == 8'h8e ? _GEN_116 : _GEN_115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_118 = ~io_inputBit | _GEN_117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_119 = i == 8'h8f ? _GEN_118 : _GEN_117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_120 = io_inputBit ? 1'h0 : _GEN_119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_121 = i == 8'h8f ? _GEN_120 : _GEN_119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_122 = ~io_inputBit ? 1'h0 : _GEN_121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_123 = i == 8'h91 ? _GEN_122 : _GEN_121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_124 = io_inputBit | _GEN_123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_125 = i == 8'h91 ? _GEN_124 : _GEN_123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_126 = ~io_inputBit | _GEN_125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_127 = i == 8'h92 ? _GEN_126 : _GEN_125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_128 = io_inputBit ? 1'h0 : _GEN_127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_129 = i == 8'h92 ? _GEN_128 : _GEN_127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_130 = io_inputBit ? 1'h0 : buffer_4; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_131 = i == 8'h0 ? _GEN_130 : buffer_4; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_132 = io_inputBit ? 1'h0 : _GEN_131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_133 = i == 8'h1 ? _GEN_132 : _GEN_131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_134 = ~io_inputBit | _GEN_133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_135 = i == 8'h7 ? _GEN_134 : _GEN_133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_136 = io_inputBit ? 1'h0 : _GEN_135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_137 = i == 8'h8 ? _GEN_136 : _GEN_135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_138 = io_inputBit ? 1'h0 : _GEN_137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_139 = i == 8'h11 ? _GEN_138 : _GEN_137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_140 = ~io_inputBit | _GEN_139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_141 = i == 8'h21 ? _GEN_140 : _GEN_139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_142 = ~io_inputBit | _GEN_141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_143 = i == 8'h44 ? _GEN_142 : _GEN_141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_144 = ~io_inputBit ? 1'h0 : _GEN_143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_145 = i == 8'h45 ? _GEN_144 : _GEN_143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_146 = ~io_inputBit | _GEN_145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_147 = i == 8'h46 ? _GEN_146 : _GEN_145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_148 = ~io_inputBit ? 1'h0 : _GEN_147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_149 = i == 8'h47 ? _GEN_148 : _GEN_147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_150 = ~io_inputBit | _GEN_149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_151 = i == 8'h48 ? _GEN_150 : _GEN_149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_152 = ~io_inputBit ? 1'h0 : _GEN_151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_153 = i == 8'h8a ? _GEN_152 : _GEN_151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_154 = io_inputBit | _GEN_153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_155 = i == 8'h8a ? _GEN_154 : _GEN_153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_156 = ~io_inputBit | _GEN_155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_157 = i == 8'h8c ? _GEN_156 : _GEN_155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_158 = io_inputBit ? 1'h0 : _GEN_157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_159 = i == 8'h8c ? _GEN_158 : _GEN_157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_160 = ~io_inputBit ? 1'h0 : _GEN_159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_161 = i == 8'h8e ? _GEN_160 : _GEN_159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_162 = io_inputBit | _GEN_161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_163 = i == 8'h8e ? _GEN_162 : _GEN_161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_164 = ~io_inputBit | _GEN_163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_165 = i == 8'h90 ? _GEN_164 : _GEN_163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_166 = io_inputBit ? 1'h0 : _GEN_165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_167 = i == 8'h90 ? _GEN_166 : _GEN_165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_168 = ~io_inputBit ? 1'h0 : _GEN_167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_169 = i == 8'h92 ? _GEN_168 : _GEN_167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_170 = io_inputBit | _GEN_169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_171 = i == 8'h92 ? _GEN_170 : _GEN_169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_172 = io_inputBit ? 1'h0 : buffer_5; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_173 = i == 8'h0 ? _GEN_172 : buffer_5; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_174 = io_inputBit ? 1'h0 : _GEN_173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_175 = i == 8'h1 ? _GEN_174 : _GEN_173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_176 = ~io_inputBit ? 1'h0 : _GEN_175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_177 = i == 8'h7 ? _GEN_176 : _GEN_175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_178 = io_inputBit ? 1'h0 : _GEN_177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_179 = i == 8'h8 ? _GEN_178 : _GEN_177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_180 = io_inputBit ? 1'h0 : _GEN_179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_181 = i == 8'h11 ? _GEN_180 : _GEN_179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_182 = ~io_inputBit ? 1'h0 : _GEN_181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_183 = i == 8'h21 ? _GEN_182 : _GEN_181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_184 = ~io_inputBit ? 1'h0 : _GEN_183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_185 = i == 8'h89 ? _GEN_184 : _GEN_183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_186 = io_inputBit | _GEN_185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_187 = i == 8'h89 ? _GEN_186 : _GEN_185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_188 = ~io_inputBit | _GEN_187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_189 = i == 8'h8a ? _GEN_188 : _GEN_187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_190 = io_inputBit ? 1'h0 : _GEN_189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_191 = i == 8'h8a ? _GEN_190 : _GEN_189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_192 = ~io_inputBit ? 1'h0 : _GEN_191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_193 = i == 8'h8b ? _GEN_192 : _GEN_191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_194 = io_inputBit | _GEN_193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_195 = i == 8'h8b ? _GEN_194 : _GEN_193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_196 = ~io_inputBit | _GEN_195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_197 = i == 8'h8c ? _GEN_196 : _GEN_195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_198 = io_inputBit ? 1'h0 : _GEN_197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_199 = i == 8'h8c ? _GEN_198 : _GEN_197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_200 = ~io_inputBit ? 1'h0 : _GEN_199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_201 = i == 8'h8d ? _GEN_200 : _GEN_199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_202 = io_inputBit | _GEN_201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_203 = i == 8'h8d ? _GEN_202 : _GEN_201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_204 = ~io_inputBit | _GEN_203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_205 = i == 8'h8e ? _GEN_204 : _GEN_203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_206 = io_inputBit ? 1'h0 : _GEN_205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_207 = i == 8'h8e ? _GEN_206 : _GEN_205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_208 = ~io_inputBit ? 1'h0 : _GEN_207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_209 = i == 8'h8f ? _GEN_208 : _GEN_207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_210 = io_inputBit | _GEN_209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_211 = i == 8'h8f ? _GEN_210 : _GEN_209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_212 = ~io_inputBit | _GEN_211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_213 = i == 8'h90 ? _GEN_212 : _GEN_211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_214 = io_inputBit ? 1'h0 : _GEN_213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_215 = i == 8'h90 ? _GEN_214 : _GEN_213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_216 = ~io_inputBit ? 1'h0 : _GEN_215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_217 = i == 8'h91 ? _GEN_216 : _GEN_215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_218 = io_inputBit | _GEN_217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_219 = i == 8'h91 ? _GEN_218 : _GEN_217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_220 = ~io_inputBit | _GEN_219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_221 = i == 8'h92 ? _GEN_220 : _GEN_219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_222 = io_inputBit ? 1'h0 : _GEN_221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_223 = i == 8'h92 ? _GEN_222 : _GEN_221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_224 = io_inputBit ? 1'h0 : buffer_6; // @[lut_mem_online.scala 209:19 236:46 238:32]
  wire  _GEN_225 = i == 8'h0 ? _GEN_224 : buffer_6; // @[lut_mem_online.scala 209:19 234:34]
  wire  _GEN_226 = io_inputBit ? 1'h0 : _GEN_225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_227 = i == 8'h1 ? _GEN_226 : _GEN_225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_228 = ~io_inputBit ? 1'h0 : _GEN_227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_229 = i == 8'h7 ? _GEN_228 : _GEN_227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_230 = io_inputBit ? 1'h0 : _GEN_229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_231 = i == 8'h8 ? _GEN_230 : _GEN_229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_232 = io_inputBit ? 1'h0 : _GEN_231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_233 = i == 8'h11 ? _GEN_232 : _GEN_231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_234 = ~io_inputBit ? 1'h0 : _GEN_233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_235 = i == 8'h21 ? _GEN_234 : _GEN_233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_236 = ~io_inputBit ? 1'h0 : _GEN_235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_237 = i == 8'h89 ? _GEN_236 : _GEN_235; // @[lut_mem_online.scala 234:34]
  wire  _GEN_238 = io_inputBit | _GEN_237; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_239 = i == 8'h89 ? _GEN_238 : _GEN_237; // @[lut_mem_online.scala 234:34]
  wire  _GEN_240 = ~io_inputBit ? 1'h0 : _GEN_239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_241 = i == 8'h8a ? _GEN_240 : _GEN_239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_242 = io_inputBit | _GEN_241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_243 = i == 8'h8a ? _GEN_242 : _GEN_241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_244 = ~io_inputBit ? 1'h0 : _GEN_243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_245 = i == 8'h8b ? _GEN_244 : _GEN_243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_246 = io_inputBit | _GEN_245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_247 = i == 8'h8b ? _GEN_246 : _GEN_245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_248 = ~io_inputBit ? 1'h0 : _GEN_247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_249 = i == 8'h8c ? _GEN_248 : _GEN_247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_250 = io_inputBit | _GEN_249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_251 = i == 8'h8c ? _GEN_250 : _GEN_249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_252 = ~io_inputBit ? 1'h0 : _GEN_251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_253 = i == 8'h8d ? _GEN_252 : _GEN_251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_254 = io_inputBit | _GEN_253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_255 = i == 8'h8d ? _GEN_254 : _GEN_253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_256 = ~io_inputBit ? 1'h0 : _GEN_255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_257 = i == 8'h8e ? _GEN_256 : _GEN_255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_258 = io_inputBit | _GEN_257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_259 = i == 8'h8e ? _GEN_258 : _GEN_257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_260 = ~io_inputBit ? 1'h0 : _GEN_259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_261 = i == 8'h8f ? _GEN_260 : _GEN_259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_262 = io_inputBit | _GEN_261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_263 = i == 8'h8f ? _GEN_262 : _GEN_261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_264 = ~io_inputBit ? 1'h0 : _GEN_263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_265 = i == 8'h90 ? _GEN_264 : _GEN_263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_266 = io_inputBit | _GEN_265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_267 = i == 8'h90 ? _GEN_266 : _GEN_265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_268 = ~io_inputBit ? 1'h0 : _GEN_267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_269 = i == 8'h91 ? _GEN_268 : _GEN_267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_270 = io_inputBit | _GEN_269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_271 = i == 8'h91 ? _GEN_270 : _GEN_269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_272 = ~io_inputBit ? 1'h0 : _GEN_271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_273 = i == 8'h92 ? _GEN_272 : _GEN_271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_274 = io_inputBit | _GEN_273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_275 = i == 8'h92 ? _GEN_274 : _GEN_273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_276 = io_inputBit ? 1'h0 : _GEN_13; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_277 = i == 8'h0 ? _GEN_276 : _GEN_13; // @[lut_mem_online.scala 234:34]
  wire  _GEN_278 = ~io_inputBit ? 1'h0 : _GEN_277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_279 = i == 8'h3 ? _GEN_278 : _GEN_277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_280 = io_inputBit ? 1'h0 : _GEN_279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_281 = i == 8'h4 ? _GEN_280 : _GEN_279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_282 = io_inputBit | _GEN_281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_283 = i == 8'h8 ? _GEN_282 : _GEN_281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_284 = io_inputBit ? 1'h0 : _GEN_283; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_285 = i == 8'h9 ? _GEN_284 : _GEN_283; // @[lut_mem_online.scala 234:34]
  wire  _GEN_286 = io_inputBit | _GEN_285; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_287 = i == 8'h11 ? _GEN_286 : _GEN_285; // @[lut_mem_online.scala 234:34]
  wire  _GEN_288 = io_inputBit ? 1'h0 : _GEN_287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_289 = i == 8'h13 ? _GEN_288 : _GEN_287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_290 = io_inputBit | _GEN_289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_291 = i == 8'h23 ? _GEN_290 : _GEN_289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_292 = ~io_inputBit | _GEN_291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_293 = i == 8'h27 ? _GEN_292 : _GEN_291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_294 = io_inputBit ? 1'h0 : _GEN_293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_295 = i == 8'h27 ? _GEN_294 : _GEN_293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_296 = io_inputBit | _GEN_295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_297 = i == 8'h47 ? _GEN_296 : _GEN_295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_298 = ~io_inputBit ? 1'h0 : _GEN_297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_299 = i == 8'h8f ? _GEN_298 : _GEN_297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_300 = io_inputBit | _GEN_299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_301 = i == 8'h8f ? _GEN_300 : _GEN_299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_302 = io_inputBit ? 1'h0 : _GEN_41; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_303 = i == 8'h0 ? _GEN_302 : _GEN_41; // @[lut_mem_online.scala 234:34]
  wire  _GEN_304 = io_inputBit ? 1'h0 : _GEN_303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_305 = i == 8'h4 ? _GEN_304 : _GEN_303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_306 = ~io_inputBit ? 1'h0 : _GEN_305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_307 = i == 8'h7 ? _GEN_306 : _GEN_305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_308 = io_inputBit ? 1'h0 : _GEN_307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_309 = i == 8'h9 ? _GEN_308 : _GEN_307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_310 = ~io_inputBit ? 1'h0 : _GEN_309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_311 = i == 8'h10 ? _GEN_310 : _GEN_309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_312 = io_inputBit | _GEN_311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_313 = i == 8'h11 ? _GEN_312 : _GEN_311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_314 = ~io_inputBit | _GEN_313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_315 = i == 8'h12 ? _GEN_314 : _GEN_313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_316 = io_inputBit | _GEN_315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_317 = i == 8'h22 ? _GEN_316 : _GEN_315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_318 = io_inputBit ? 1'h0 : _GEN_317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_319 = i == 8'h23 ? _GEN_318 : _GEN_317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_320 = ~io_inputBit | _GEN_319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_321 = i == 8'h26 ? _GEN_320 : _GEN_319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_322 = ~io_inputBit ? 1'h0 : _GEN_321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_323 = i == 8'h27 ? _GEN_322 : _GEN_321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_324 = io_inputBit | _GEN_323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_325 = i == 8'h27 ? _GEN_324 : _GEN_323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_326 = io_inputBit ? 1'h0 : _GEN_325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_327 = i == 8'h28 ? _GEN_326 : _GEN_325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_328 = ~io_inputBit ? 1'h0 : _GEN_327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_329 = i == 8'h45 ? _GEN_328 : _GEN_327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_330 = io_inputBit ? 1'h0 : _GEN_329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_331 = i == 8'h47 ? _GEN_330 : _GEN_329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_332 = io_inputBit ? 1'h0 : _GEN_331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_333 = i == 8'h4e ? _GEN_332 : _GEN_331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_334 = ~io_inputBit | _GEN_333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_335 = i == 8'h51 ? _GEN_334 : _GEN_333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_336 = io_inputBit ? 1'h0 : _GEN_335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_337 = i == 8'h51 ? _GEN_336 : _GEN_335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_338 = ~io_inputBit ? 1'h0 : _GEN_337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_339 = i == 8'h8c ? _GEN_338 : _GEN_337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_340 = io_inputBit | _GEN_339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_341 = i == 8'h8c ? _GEN_340 : _GEN_339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_342 = ~io_inputBit | _GEN_341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_343 = i == 8'h8f ? _GEN_342 : _GEN_341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_344 = io_inputBit ? 1'h0 : _GEN_343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_345 = i == 8'h8f ? _GEN_344 : _GEN_343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_346 = ~io_inputBit | _GEN_345; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_347 = i == 8'h9d ? _GEN_346 : _GEN_345; // @[lut_mem_online.scala 234:34]
  wire  _GEN_348 = io_inputBit ? 1'h0 : _GEN_347; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_349 = i == 8'h9d ? _GEN_348 : _GEN_347; // @[lut_mem_online.scala 234:34]
  wire  _GEN_350 = io_inputBit ? 1'h0 : _GEN_81; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_351 = i == 8'h0 ? _GEN_350 : _GEN_81; // @[lut_mem_online.scala 234:34]
  wire  _GEN_352 = io_inputBit ? 1'h0 : _GEN_351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_353 = i == 8'h4 ? _GEN_352 : _GEN_351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_354 = ~io_inputBit ? 1'h0 : _GEN_353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_355 = i == 8'h7 ? _GEN_354 : _GEN_353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_356 = io_inputBit ? 1'h0 : _GEN_355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_357 = i == 8'h9 ? _GEN_356 : _GEN_355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_358 = ~io_inputBit ? 1'h0 : _GEN_357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_359 = i == 8'h10 ? _GEN_358 : _GEN_357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_360 = io_inputBit ? 1'h0 : _GEN_359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_361 = i == 8'h11 ? _GEN_360 : _GEN_359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_362 = ~io_inputBit ? 1'h0 : _GEN_361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_363 = i == 8'h12 ? _GEN_362 : _GEN_361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_364 = io_inputBit | _GEN_363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_365 = i == 8'h23 ? _GEN_364 : _GEN_363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_366 = ~io_inputBit ? 1'h0 : _GEN_365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_367 = i == 8'h26 ? _GEN_366 : _GEN_365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_368 = ~io_inputBit | _GEN_367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_369 = i == 8'h45 ? _GEN_368 : _GEN_367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_370 = ~io_inputBit ? 1'h0 : _GEN_369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_371 = i == 8'h46 ? _GEN_370 : _GEN_369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_372 = io_inputBit | _GEN_371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_373 = i == 8'h46 ? _GEN_372 : _GEN_371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_374 = io_inputBit ? 1'h0 : _GEN_373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_375 = i == 8'h47 ? _GEN_374 : _GEN_373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_376 = io_inputBit | _GEN_375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_377 = i == 8'h4e ? _GEN_376 : _GEN_375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_378 = io_inputBit ? 1'h0 : _GEN_377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_379 = i == 8'h4f ? _GEN_378 : _GEN_377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_380 = ~io_inputBit | _GEN_379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_381 = i == 8'h50 ? _GEN_380 : _GEN_379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_382 = ~io_inputBit ? 1'h0 : _GEN_381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_383 = i == 8'h51 ? _GEN_382 : _GEN_381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_384 = io_inputBit | _GEN_383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_385 = i == 8'h51 ? _GEN_384 : _GEN_383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_386 = io_inputBit ? 1'h0 : _GEN_385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_387 = i == 8'h52 ? _GEN_386 : _GEN_385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_388 = ~io_inputBit | _GEN_387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_389 = i == 8'h8c ? _GEN_388 : _GEN_387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_390 = io_inputBit ? 1'h0 : _GEN_389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_391 = i == 8'h8c ? _GEN_390 : _GEN_389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_392 = ~io_inputBit | _GEN_391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_393 = i == 8'h8f ? _GEN_392 : _GEN_391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_394 = io_inputBit ? 1'h0 : _GEN_393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_395 = i == 8'h8f ? _GEN_394 : _GEN_393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_396 = ~io_inputBit ? 1'h0 : _GEN_395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_397 = i == 8'h9d ? _GEN_396 : _GEN_395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_398 = io_inputBit | _GEN_397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_399 = i == 8'h9d ? _GEN_398 : _GEN_397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_400 = ~io_inputBit | _GEN_399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_401 = i == 8'h9f ? _GEN_400 : _GEN_399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_402 = io_inputBit ? 1'h0 : _GEN_401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_403 = i == 8'h9f ? _GEN_402 : _GEN_401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_404 = ~io_inputBit | _GEN_403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_405 = i == 8'ha2 ? _GEN_404 : _GEN_403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_406 = io_inputBit ? 1'h0 : _GEN_405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_407 = i == 8'ha2 ? _GEN_406 : _GEN_405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_408 = ~io_inputBit | _GEN_407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_409 = i == 8'ha5 ? _GEN_408 : _GEN_407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_410 = io_inputBit ? 1'h0 : _GEN_409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_411 = i == 8'ha5 ? _GEN_410 : _GEN_409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_412 = io_inputBit ? 1'h0 : _GEN_129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_413 = i == 8'h0 ? _GEN_412 : _GEN_129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_414 = io_inputBit ? 1'h0 : _GEN_413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_415 = i == 8'h4 ? _GEN_414 : _GEN_413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_416 = ~io_inputBit ? 1'h0 : _GEN_415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_417 = i == 8'h7 ? _GEN_416 : _GEN_415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_418 = io_inputBit ? 1'h0 : _GEN_417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_419 = i == 8'h9 ? _GEN_418 : _GEN_417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_420 = io_inputBit ? 1'h0 : _GEN_419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_421 = i == 8'h11 ? _GEN_420 : _GEN_419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_422 = ~io_inputBit ? 1'h0 : _GEN_421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_423 = i == 8'h12 ? _GEN_422 : _GEN_421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_424 = ~io_inputBit ? 1'h0 : _GEN_423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_425 = i == 8'h21 ? _GEN_424 : _GEN_423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_426 = ~io_inputBit ? 1'h0 : _GEN_425; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_427 = i == 8'h26 ? _GEN_426 : _GEN_425; // @[lut_mem_online.scala 234:34]
  wire  _GEN_428 = ~io_inputBit ? 1'h0 : _GEN_427; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_429 = i == 8'h44 ? _GEN_428 : _GEN_427; // @[lut_mem_online.scala 234:34]
  wire  _GEN_430 = io_inputBit | _GEN_429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_431 = i == 8'h44 ? _GEN_430 : _GEN_429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_432 = ~io_inputBit | _GEN_431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_433 = i == 8'h46 ? _GEN_432 : _GEN_431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_434 = io_inputBit ? 1'h0 : _GEN_433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_435 = i == 8'h46 ? _GEN_434 : _GEN_433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_436 = ~io_inputBit ? 1'h0 : _GEN_435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_437 = i == 8'h48 ? _GEN_436 : _GEN_435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_438 = io_inputBit | _GEN_437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_439 = i == 8'h48 ? _GEN_438 : _GEN_437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_440 = io_inputBit ? 1'h0 : _GEN_439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_441 = i == 8'h4f ? _GEN_440 : _GEN_439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_442 = io_inputBit | _GEN_441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_443 = i == 8'h51 ? _GEN_442 : _GEN_441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_444 = ~io_inputBit ? 1'h0 : _GEN_443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_445 = i == 8'h8b ? _GEN_444 : _GEN_443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_446 = io_inputBit | _GEN_445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_447 = i == 8'h8b ? _GEN_446 : _GEN_445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_448 = ~io_inputBit | _GEN_447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_449 = i == 8'h8c ? _GEN_448 : _GEN_447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_450 = io_inputBit ? 1'h0 : _GEN_449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_451 = i == 8'h8c ? _GEN_450 : _GEN_449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_452 = ~io_inputBit | _GEN_451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_453 = i == 8'h8f ? _GEN_452 : _GEN_451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_454 = io_inputBit ? 1'h0 : _GEN_453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_455 = i == 8'h8f ? _GEN_454 : _GEN_453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_456 = ~io_inputBit ? 1'h0 : _GEN_455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_457 = i == 8'h90 ? _GEN_456 : _GEN_455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_458 = io_inputBit | _GEN_457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_459 = i == 8'h90 ? _GEN_458 : _GEN_457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_460 = ~io_inputBit ? 1'h0 : _GEN_459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_461 = i == 8'h9d ? _GEN_460 : _GEN_459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_462 = io_inputBit | _GEN_461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_463 = i == 8'h9d ? _GEN_462 : _GEN_461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_464 = ~io_inputBit | _GEN_463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_465 = i == 8'h9e ? _GEN_464 : _GEN_463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_466 = io_inputBit ? 1'h0 : _GEN_465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_467 = i == 8'h9e ? _GEN_466 : _GEN_465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_468 = ~io_inputBit ? 1'h0 : _GEN_467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_469 = i == 8'h9f ? _GEN_468 : _GEN_467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_470 = io_inputBit | _GEN_469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_471 = i == 8'h9f ? _GEN_470 : _GEN_469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_472 = ~io_inputBit | _GEN_471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_473 = i == 8'ha1 ? _GEN_472 : _GEN_471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_474 = io_inputBit ? 1'h0 : _GEN_473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_475 = i == 8'ha1 ? _GEN_474 : _GEN_473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_476 = ~io_inputBit ? 1'h0 : _GEN_475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_477 = i == 8'ha2 ? _GEN_476 : _GEN_475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_478 = io_inputBit | _GEN_477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_479 = i == 8'ha2 ? _GEN_478 : _GEN_477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_480 = ~io_inputBit | _GEN_479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_481 = i == 8'ha3 ? _GEN_480 : _GEN_479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_482 = io_inputBit ? 1'h0 : _GEN_481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_483 = i == 8'ha3 ? _GEN_482 : _GEN_481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_484 = ~io_inputBit ? 1'h0 : _GEN_483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_485 = i == 8'ha5 ? _GEN_484 : _GEN_483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_486 = io_inputBit | _GEN_485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_487 = i == 8'ha5 ? _GEN_486 : _GEN_485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_488 = ~io_inputBit | _GEN_487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_489 = i == 8'ha6 ? _GEN_488 : _GEN_487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_490 = io_inputBit ? 1'h0 : _GEN_489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_491 = i == 8'ha6 ? _GEN_490 : _GEN_489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_492 = io_inputBit ? 1'h0 : _GEN_171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_493 = i == 8'h0 ? _GEN_492 : _GEN_171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_494 = io_inputBit ? 1'h0 : _GEN_493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_495 = i == 8'h4 ? _GEN_494 : _GEN_493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_496 = ~io_inputBit ? 1'h0 : _GEN_495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_497 = i == 8'h7 ? _GEN_496 : _GEN_495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_498 = io_inputBit ? 1'h0 : _GEN_497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_499 = i == 8'h9 ? _GEN_498 : _GEN_497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_500 = io_inputBit | _GEN_499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_501 = i == 8'h11 ? _GEN_500 : _GEN_499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_502 = ~io_inputBit | _GEN_501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_503 = i == 8'h12 ? _GEN_502 : _GEN_501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_504 = ~io_inputBit ? 1'h0 : _GEN_503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_505 = i == 8'h21 ? _GEN_504 : _GEN_503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_506 = ~io_inputBit | _GEN_505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_507 = i == 8'h26 ? _GEN_506 : _GEN_505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_508 = ~io_inputBit | _GEN_507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_509 = i == 8'h4e ? _GEN_508 : _GEN_507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_510 = ~io_inputBit ? 1'h0 : _GEN_509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_511 = i == 8'h4f ? _GEN_510 : _GEN_509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_512 = ~io_inputBit | _GEN_511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_513 = i == 8'h50 ? _GEN_512 : _GEN_511; // @[lut_mem_online.scala 234:34]
  wire  _GEN_514 = ~io_inputBit ? 1'h0 : _GEN_513; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_515 = i == 8'h51 ? _GEN_514 : _GEN_513; // @[lut_mem_online.scala 234:34]
  wire  _GEN_516 = ~io_inputBit | _GEN_515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_517 = i == 8'h52 ? _GEN_516 : _GEN_515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_518 = ~io_inputBit ? 1'h0 : _GEN_517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_519 = i == 8'h89 ? _GEN_518 : _GEN_517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_520 = io_inputBit | _GEN_519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_521 = i == 8'h89 ? _GEN_520 : _GEN_519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_522 = ~io_inputBit ? 1'h0 : _GEN_521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_523 = i == 8'h8a ? _GEN_522 : _GEN_521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_524 = io_inputBit | _GEN_523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_525 = i == 8'h8a ? _GEN_524 : _GEN_523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_526 = ~io_inputBit | _GEN_525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_527 = i == 8'h8b ? _GEN_526 : _GEN_525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_528 = io_inputBit ? 1'h0 : _GEN_527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_529 = i == 8'h8b ? _GEN_528 : _GEN_527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_530 = ~io_inputBit | _GEN_529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_531 = i == 8'h8c ? _GEN_530 : _GEN_529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_532 = io_inputBit ? 1'h0 : _GEN_531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_533 = i == 8'h8c ? _GEN_532 : _GEN_531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_534 = ~io_inputBit ? 1'h0 : _GEN_533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_535 = i == 8'h8d ? _GEN_534 : _GEN_533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_536 = io_inputBit | _GEN_535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_537 = i == 8'h8d ? _GEN_536 : _GEN_535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_538 = ~io_inputBit ? 1'h0 : _GEN_537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_539 = i == 8'h8e ? _GEN_538 : _GEN_537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_540 = io_inputBit | _GEN_539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_541 = i == 8'h8e ? _GEN_540 : _GEN_539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_542 = ~io_inputBit | _GEN_541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_543 = i == 8'h8f ? _GEN_542 : _GEN_541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_544 = io_inputBit ? 1'h0 : _GEN_543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_545 = i == 8'h8f ? _GEN_544 : _GEN_543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_546 = ~io_inputBit | _GEN_545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_547 = i == 8'h90 ? _GEN_546 : _GEN_545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_548 = io_inputBit ? 1'h0 : _GEN_547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_549 = i == 8'h90 ? _GEN_548 : _GEN_547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_550 = ~io_inputBit ? 1'h0 : _GEN_549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_551 = i == 8'h91 ? _GEN_550 : _GEN_549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_552 = io_inputBit | _GEN_551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_553 = i == 8'h91 ? _GEN_552 : _GEN_551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_554 = ~io_inputBit ? 1'h0 : _GEN_553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_555 = i == 8'h92 ? _GEN_554 : _GEN_553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_556 = io_inputBit | _GEN_555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_557 = i == 8'h92 ? _GEN_556 : _GEN_555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_558 = ~io_inputBit ? 1'h0 : _GEN_557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_559 = i == 8'h9e ? _GEN_558 : _GEN_557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_560 = io_inputBit | _GEN_559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_561 = i == 8'h9e ? _GEN_560 : _GEN_559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_562 = ~io_inputBit | _GEN_561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_563 = i == 8'ha0 ? _GEN_562 : _GEN_561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_564 = io_inputBit ? 1'h0 : _GEN_563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_565 = i == 8'ha0 ? _GEN_564 : _GEN_563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_566 = ~io_inputBit ? 1'h0 : _GEN_565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_567 = i == 8'ha2 ? _GEN_566 : _GEN_565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_568 = io_inputBit | _GEN_567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_569 = i == 8'ha2 ? _GEN_568 : _GEN_567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_570 = ~io_inputBit | _GEN_569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_571 = i == 8'ha4 ? _GEN_570 : _GEN_569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_572 = io_inputBit ? 1'h0 : _GEN_571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_573 = i == 8'ha4 ? _GEN_572 : _GEN_571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_574 = ~io_inputBit ? 1'h0 : _GEN_573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_575 = i == 8'ha6 ? _GEN_574 : _GEN_573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_576 = io_inputBit | _GEN_575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_577 = i == 8'ha6 ? _GEN_576 : _GEN_575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_578 = io_inputBit ? 1'h0 : _GEN_223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_579 = i == 8'h0 ? _GEN_578 : _GEN_223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_580 = io_inputBit ? 1'h0 : _GEN_579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_581 = i == 8'h4 ? _GEN_580 : _GEN_579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_582 = ~io_inputBit ? 1'h0 : _GEN_581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_583 = i == 8'h7 ? _GEN_582 : _GEN_581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_584 = io_inputBit ? 1'h0 : _GEN_583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_585 = i == 8'h9 ? _GEN_584 : _GEN_583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_586 = io_inputBit ? 1'h0 : _GEN_585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_587 = i == 8'h11 ? _GEN_586 : _GEN_585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_588 = ~io_inputBit ? 1'h0 : _GEN_587; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_589 = i == 8'h12 ? _GEN_588 : _GEN_587; // @[lut_mem_online.scala 234:34]
  wire  _GEN_590 = ~io_inputBit ? 1'h0 : _GEN_589; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_591 = i == 8'h21 ? _GEN_590 : _GEN_589; // @[lut_mem_online.scala 234:34]
  wire  _GEN_592 = ~io_inputBit ? 1'h0 : _GEN_591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_593 = i == 8'h26 ? _GEN_592 : _GEN_591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_594 = ~io_inputBit ? 1'h0 : _GEN_593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_595 = i == 8'h44 ? _GEN_594 : _GEN_593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_596 = io_inputBit | _GEN_595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_597 = i == 8'h44 ? _GEN_596 : _GEN_595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_598 = ~io_inputBit ? 1'h0 : _GEN_597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_599 = i == 8'h45 ? _GEN_598 : _GEN_597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_600 = io_inputBit | _GEN_599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_601 = i == 8'h45 ? _GEN_600 : _GEN_599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_602 = ~io_inputBit ? 1'h0 : _GEN_601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_603 = i == 8'h46 ? _GEN_602 : _GEN_601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_604 = io_inputBit | _GEN_603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_605 = i == 8'h46 ? _GEN_604 : _GEN_603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_606 = ~io_inputBit ? 1'h0 : _GEN_605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_607 = i == 8'h47 ? _GEN_606 : _GEN_605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_608 = io_inputBit | _GEN_607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_609 = i == 8'h47 ? _GEN_608 : _GEN_607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_610 = ~io_inputBit ? 1'h0 : _GEN_609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_611 = i == 8'h48 ? _GEN_610 : _GEN_609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_612 = io_inputBit | _GEN_611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_613 = i == 8'h48 ? _GEN_612 : _GEN_611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_614 = ~io_inputBit ? 1'h0 : _GEN_613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_615 = i == 8'h9d ? _GEN_614 : _GEN_613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_616 = io_inputBit | _GEN_615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_617 = i == 8'h9d ? _GEN_616 : _GEN_615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_618 = ~io_inputBit | _GEN_617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_619 = i == 8'h9e ? _GEN_618 : _GEN_617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_620 = io_inputBit ? 1'h0 : _GEN_619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_621 = i == 8'h9e ? _GEN_620 : _GEN_619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_622 = ~io_inputBit ? 1'h0 : _GEN_621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_623 = i == 8'h9f ? _GEN_622 : _GEN_621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_624 = io_inputBit | _GEN_623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_625 = i == 8'h9f ? _GEN_624 : _GEN_623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_626 = ~io_inputBit | _GEN_625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_627 = i == 8'ha0 ? _GEN_626 : _GEN_625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_628 = io_inputBit ? 1'h0 : _GEN_627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_629 = i == 8'ha0 ? _GEN_628 : _GEN_627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_630 = ~io_inputBit ? 1'h0 : _GEN_629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_631 = i == 8'ha1 ? _GEN_630 : _GEN_629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_632 = io_inputBit | _GEN_631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_633 = i == 8'ha1 ? _GEN_632 : _GEN_631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_634 = ~io_inputBit | _GEN_633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_635 = i == 8'ha2 ? _GEN_634 : _GEN_633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_636 = io_inputBit ? 1'h0 : _GEN_635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_637 = i == 8'ha2 ? _GEN_636 : _GEN_635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_638 = ~io_inputBit ? 1'h0 : _GEN_637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_639 = i == 8'ha3 ? _GEN_638 : _GEN_637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_640 = io_inputBit | _GEN_639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_641 = i == 8'ha3 ? _GEN_640 : _GEN_639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_642 = ~io_inputBit | _GEN_641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_643 = i == 8'ha4 ? _GEN_642 : _GEN_641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_644 = io_inputBit ? 1'h0 : _GEN_643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_645 = i == 8'ha4 ? _GEN_644 : _GEN_643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_646 = ~io_inputBit ? 1'h0 : _GEN_645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_647 = i == 8'ha5 ? _GEN_646 : _GEN_645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_648 = io_inputBit | _GEN_647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_649 = i == 8'ha5 ? _GEN_648 : _GEN_647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_650 = ~io_inputBit | _GEN_649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_651 = i == 8'ha6 ? _GEN_650 : _GEN_649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_652 = io_inputBit ? 1'h0 : _GEN_651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_653 = i == 8'ha6 ? _GEN_652 : _GEN_651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_654 = io_inputBit ? 1'h0 : _GEN_275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_655 = i == 8'h0 ? _GEN_654 : _GEN_275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_656 = io_inputBit ? 1'h0 : _GEN_655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_657 = i == 8'h4 ? _GEN_656 : _GEN_655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_658 = ~io_inputBit ? 1'h0 : _GEN_657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_659 = i == 8'h7 ? _GEN_658 : _GEN_657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_660 = io_inputBit ? 1'h0 : _GEN_659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_661 = i == 8'h9 ? _GEN_660 : _GEN_659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_662 = io_inputBit ? 1'h0 : _GEN_661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_663 = i == 8'h11 ? _GEN_662 : _GEN_661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_664 = ~io_inputBit ? 1'h0 : _GEN_663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_665 = i == 8'h12 ? _GEN_664 : _GEN_663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_666 = ~io_inputBit ? 1'h0 : _GEN_665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_667 = i == 8'h21 ? _GEN_666 : _GEN_665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_668 = ~io_inputBit ? 1'h0 : _GEN_667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_669 = i == 8'h26 ? _GEN_668 : _GEN_667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_670 = ~io_inputBit ? 1'h0 : _GEN_669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_671 = i == 8'h89 ? _GEN_670 : _GEN_669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_672 = io_inputBit | _GEN_671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_673 = i == 8'h89 ? _GEN_672 : _GEN_671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_674 = ~io_inputBit ? 1'h0 : _GEN_673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_675 = i == 8'h8a ? _GEN_674 : _GEN_673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_676 = io_inputBit | _GEN_675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_677 = i == 8'h8a ? _GEN_676 : _GEN_675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_678 = ~io_inputBit ? 1'h0 : _GEN_677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_679 = i == 8'h8b ? _GEN_678 : _GEN_677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_680 = io_inputBit | _GEN_679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_681 = i == 8'h8b ? _GEN_680 : _GEN_679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_682 = ~io_inputBit ? 1'h0 : _GEN_681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_683 = i == 8'h8c ? _GEN_682 : _GEN_681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_684 = io_inputBit | _GEN_683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_685 = i == 8'h8c ? _GEN_684 : _GEN_683; // @[lut_mem_online.scala 234:34]
  wire  _GEN_686 = ~io_inputBit ? 1'h0 : _GEN_685; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_687 = i == 8'h8d ? _GEN_686 : _GEN_685; // @[lut_mem_online.scala 234:34]
  wire  _GEN_688 = io_inputBit | _GEN_687; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_689 = i == 8'h8d ? _GEN_688 : _GEN_687; // @[lut_mem_online.scala 234:34]
  wire  _GEN_690 = ~io_inputBit ? 1'h0 : _GEN_689; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_691 = i == 8'h8e ? _GEN_690 : _GEN_689; // @[lut_mem_online.scala 234:34]
  wire  _GEN_692 = io_inputBit | _GEN_691; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_693 = i == 8'h8e ? _GEN_692 : _GEN_691; // @[lut_mem_online.scala 234:34]
  wire  _GEN_694 = ~io_inputBit ? 1'h0 : _GEN_693; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_695 = i == 8'h8f ? _GEN_694 : _GEN_693; // @[lut_mem_online.scala 234:34]
  wire  _GEN_696 = io_inputBit | _GEN_695; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_697 = i == 8'h8f ? _GEN_696 : _GEN_695; // @[lut_mem_online.scala 234:34]
  wire  _GEN_698 = ~io_inputBit ? 1'h0 : _GEN_697; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_699 = i == 8'h90 ? _GEN_698 : _GEN_697; // @[lut_mem_online.scala 234:34]
  wire  _GEN_700 = io_inputBit | _GEN_699; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_701 = i == 8'h90 ? _GEN_700 : _GEN_699; // @[lut_mem_online.scala 234:34]
  wire  _GEN_702 = ~io_inputBit ? 1'h0 : _GEN_701; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_703 = i == 8'h91 ? _GEN_702 : _GEN_701; // @[lut_mem_online.scala 234:34]
  wire  _GEN_704 = io_inputBit | _GEN_703; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_705 = i == 8'h91 ? _GEN_704 : _GEN_703; // @[lut_mem_online.scala 234:34]
  wire  _GEN_706 = ~io_inputBit ? 1'h0 : _GEN_705; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_707 = i == 8'h92 ? _GEN_706 : _GEN_705; // @[lut_mem_online.scala 234:34]
  wire  _GEN_708 = io_inputBit | _GEN_707; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_709 = i == 8'h92 ? _GEN_708 : _GEN_707; // @[lut_mem_online.scala 234:34]
  wire  _GEN_710 = ~io_inputBit ? 1'h0 : _GEN_709; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_711 = i == 8'h9d ? _GEN_710 : _GEN_709; // @[lut_mem_online.scala 234:34]
  wire  _GEN_712 = io_inputBit | _GEN_711; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_713 = i == 8'h9d ? _GEN_712 : _GEN_711; // @[lut_mem_online.scala 234:34]
  wire  _GEN_714 = ~io_inputBit ? 1'h0 : _GEN_713; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_715 = i == 8'h9e ? _GEN_714 : _GEN_713; // @[lut_mem_online.scala 234:34]
  wire  _GEN_716 = io_inputBit | _GEN_715; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_717 = i == 8'h9e ? _GEN_716 : _GEN_715; // @[lut_mem_online.scala 234:34]
  wire  _GEN_718 = ~io_inputBit ? 1'h0 : _GEN_717; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_719 = i == 8'h9f ? _GEN_718 : _GEN_717; // @[lut_mem_online.scala 234:34]
  wire  _GEN_720 = io_inputBit | _GEN_719; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_721 = i == 8'h9f ? _GEN_720 : _GEN_719; // @[lut_mem_online.scala 234:34]
  wire  _GEN_722 = ~io_inputBit ? 1'h0 : _GEN_721; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_723 = i == 8'ha0 ? _GEN_722 : _GEN_721; // @[lut_mem_online.scala 234:34]
  wire  _GEN_724 = io_inputBit | _GEN_723; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_725 = i == 8'ha0 ? _GEN_724 : _GEN_723; // @[lut_mem_online.scala 234:34]
  wire  _GEN_726 = ~io_inputBit ? 1'h0 : _GEN_725; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_727 = i == 8'ha1 ? _GEN_726 : _GEN_725; // @[lut_mem_online.scala 234:34]
  wire  _GEN_728 = io_inputBit | _GEN_727; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_729 = i == 8'ha1 ? _GEN_728 : _GEN_727; // @[lut_mem_online.scala 234:34]
  wire  _GEN_730 = ~io_inputBit ? 1'h0 : _GEN_729; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_731 = i == 8'ha2 ? _GEN_730 : _GEN_729; // @[lut_mem_online.scala 234:34]
  wire  _GEN_732 = io_inputBit | _GEN_731; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_733 = i == 8'ha2 ? _GEN_732 : _GEN_731; // @[lut_mem_online.scala 234:34]
  wire  _GEN_734 = ~io_inputBit ? 1'h0 : _GEN_733; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_735 = i == 8'ha3 ? _GEN_734 : _GEN_733; // @[lut_mem_online.scala 234:34]
  wire  _GEN_736 = io_inputBit | _GEN_735; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_737 = i == 8'ha3 ? _GEN_736 : _GEN_735; // @[lut_mem_online.scala 234:34]
  wire  _GEN_738 = ~io_inputBit ? 1'h0 : _GEN_737; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_739 = i == 8'ha4 ? _GEN_738 : _GEN_737; // @[lut_mem_online.scala 234:34]
  wire  _GEN_740 = io_inputBit | _GEN_739; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_741 = i == 8'ha4 ? _GEN_740 : _GEN_739; // @[lut_mem_online.scala 234:34]
  wire  _GEN_742 = ~io_inputBit ? 1'h0 : _GEN_741; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_743 = i == 8'ha5 ? _GEN_742 : _GEN_741; // @[lut_mem_online.scala 234:34]
  wire  _GEN_744 = io_inputBit | _GEN_743; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_745 = i == 8'ha5 ? _GEN_744 : _GEN_743; // @[lut_mem_online.scala 234:34]
  wire  _GEN_746 = ~io_inputBit ? 1'h0 : _GEN_745; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_747 = i == 8'ha6 ? _GEN_746 : _GEN_745; // @[lut_mem_online.scala 234:34]
  wire  _GEN_748 = io_inputBit | _GEN_747; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_749 = i == 8'ha6 ? _GEN_748 : _GEN_747; // @[lut_mem_online.scala 234:34]
  wire  _GEN_750 = io_inputBit ? 1'h0 : _GEN_301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_751 = i == 8'h0 ? _GEN_750 : _GEN_301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_752 = ~io_inputBit ? 1'h0 : _GEN_751; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_753 = i == 8'h1 ? _GEN_752 : _GEN_751; // @[lut_mem_online.scala 234:34]
  wire  _GEN_754 = io_inputBit | _GEN_753; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_755 = i == 8'h9 ? _GEN_754 : _GEN_753; // @[lut_mem_online.scala 234:34]
  wire  _GEN_756 = io_inputBit ? 1'h0 : _GEN_755; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_757 = i == 8'ha ? _GEN_756 : _GEN_755; // @[lut_mem_online.scala 234:34]
  wire  _GEN_758 = ~io_inputBit ? 1'h0 : _GEN_757; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_759 = i == 8'h13 ? _GEN_758 : _GEN_757; // @[lut_mem_online.scala 234:34]
  wire  _GEN_760 = ~io_inputBit | _GEN_759; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_761 = i == 8'h15 ? _GEN_760 : _GEN_759; // @[lut_mem_online.scala 234:34]
  wire  _GEN_762 = io_inputBit | _GEN_761; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_763 = i == 8'h28 ? _GEN_762 : _GEN_761; // @[lut_mem_online.scala 234:34]
  wire  _GEN_764 = ~io_inputBit | _GEN_763; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_765 = i == 8'h2c ? _GEN_764 : _GEN_763; // @[lut_mem_online.scala 234:34]
  wire  _GEN_766 = io_inputBit ? 1'h0 : _GEN_765; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_767 = i == 8'h2c ? _GEN_766 : _GEN_765; // @[lut_mem_online.scala 234:34]
  wire  _GEN_768 = io_inputBit | _GEN_767; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_769 = i == 8'h51 ? _GEN_768 : _GEN_767; // @[lut_mem_online.scala 234:34]
  wire  _GEN_770 = ~io_inputBit ? 1'h0 : _GEN_769; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_771 = i == 8'ha3 ? _GEN_770 : _GEN_769; // @[lut_mem_online.scala 234:34]
  wire  _GEN_772 = io_inputBit | _GEN_771; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_773 = i == 8'ha3 ? _GEN_772 : _GEN_771; // @[lut_mem_online.scala 234:34]
  wire  _GEN_774 = io_inputBit ? 1'h0 : _GEN_349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_775 = i == 8'h0 ? _GEN_774 : _GEN_349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_776 = ~io_inputBit ? 1'h0 : _GEN_775; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_777 = i == 8'h1 ? _GEN_776 : _GEN_775; // @[lut_mem_online.scala 234:34]
  wire  _GEN_778 = io_inputBit | _GEN_777; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_779 = i == 8'h9 ? _GEN_778 : _GEN_777; // @[lut_mem_online.scala 234:34]
  wire  _GEN_780 = io_inputBit ? 1'h0 : _GEN_779; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_781 = i == 8'h16 ? _GEN_780 : _GEN_779; // @[lut_mem_online.scala 234:34]
  wire  _GEN_782 = io_inputBit | _GEN_781; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_783 = i == 8'h27 ? _GEN_782 : _GEN_781; // @[lut_mem_online.scala 234:34]
  wire  _GEN_784 = io_inputBit ? 1'h0 : _GEN_783; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_785 = i == 8'h28 ? _GEN_784 : _GEN_783; // @[lut_mem_online.scala 234:34]
  wire  _GEN_786 = ~io_inputBit | _GEN_785; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_787 = i == 8'h2b ? _GEN_786 : _GEN_785; // @[lut_mem_online.scala 234:34]
  wire  _GEN_788 = ~io_inputBit ? 1'h0 : _GEN_787; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_789 = i == 8'h2c ? _GEN_788 : _GEN_787; // @[lut_mem_online.scala 234:34]
  wire  _GEN_790 = io_inputBit | _GEN_789; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_791 = i == 8'h2c ? _GEN_790 : _GEN_789; // @[lut_mem_online.scala 234:34]
  wire  _GEN_792 = io_inputBit ? 1'h0 : _GEN_791; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_793 = i == 8'h2d ? _GEN_792 : _GEN_791; // @[lut_mem_online.scala 234:34]
  wire  _GEN_794 = ~io_inputBit ? 1'h0 : _GEN_793; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_795 = i == 8'h4f ? _GEN_794 : _GEN_793; // @[lut_mem_online.scala 234:34]
  wire  _GEN_796 = io_inputBit ? 1'h0 : _GEN_795; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_797 = i == 8'h51 ? _GEN_796 : _GEN_795; // @[lut_mem_online.scala 234:34]
  wire  _GEN_798 = io_inputBit ? 1'h0 : _GEN_797; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_799 = i == 8'h58 ? _GEN_798 : _GEN_797; // @[lut_mem_online.scala 234:34]
  wire  _GEN_800 = ~io_inputBit | _GEN_799; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_801 = i == 8'h5b ? _GEN_800 : _GEN_799; // @[lut_mem_online.scala 234:34]
  wire  _GEN_802 = io_inputBit ? 1'h0 : _GEN_801; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_803 = i == 8'h5b ? _GEN_802 : _GEN_801; // @[lut_mem_online.scala 234:34]
  wire  _GEN_804 = ~io_inputBit ? 1'h0 : _GEN_803; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_805 = i == 8'ha0 ? _GEN_804 : _GEN_803; // @[lut_mem_online.scala 234:34]
  wire  _GEN_806 = io_inputBit | _GEN_805; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_807 = i == 8'ha0 ? _GEN_806 : _GEN_805; // @[lut_mem_online.scala 234:34]
  wire  _GEN_808 = ~io_inputBit | _GEN_807; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_809 = i == 8'ha3 ? _GEN_808 : _GEN_807; // @[lut_mem_online.scala 234:34]
  wire  _GEN_810 = io_inputBit ? 1'h0 : _GEN_809; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_811 = i == 8'ha3 ? _GEN_810 : _GEN_809; // @[lut_mem_online.scala 234:34]
  wire  _GEN_812 = ~io_inputBit | _GEN_811; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_813 = i == 8'hb1 ? _GEN_812 : _GEN_811; // @[lut_mem_online.scala 234:34]
  wire  _GEN_814 = io_inputBit ? 1'h0 : _GEN_813; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_815 = i == 8'hb1 ? _GEN_814 : _GEN_813; // @[lut_mem_online.scala 234:34]
  wire  _GEN_816 = io_inputBit ? 1'h0 : _GEN_411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_817 = i == 8'h0 ? _GEN_816 : _GEN_411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_818 = ~io_inputBit ? 1'h0 : _GEN_817; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_819 = i == 8'h1 ? _GEN_818 : _GEN_817; // @[lut_mem_online.scala 234:34]
  wire  _GEN_820 = io_inputBit ? 1'h0 : _GEN_819; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_821 = i == 8'h9 ? _GEN_820 : _GEN_819; // @[lut_mem_online.scala 234:34]
  wire  _GEN_822 = io_inputBit ? 1'h0 : _GEN_821; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_823 = i == 8'h16 ? _GEN_822 : _GEN_821; // @[lut_mem_online.scala 234:34]
  wire  _GEN_824 = io_inputBit | _GEN_823; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_825 = i == 8'h28 ? _GEN_824 : _GEN_823; // @[lut_mem_online.scala 234:34]
  wire  _GEN_826 = ~io_inputBit ? 1'h0 : _GEN_825; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_827 = i == 8'h2b ? _GEN_826 : _GEN_825; // @[lut_mem_online.scala 234:34]
  wire  _GEN_828 = ~io_inputBit | _GEN_827; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_829 = i == 8'h4f ? _GEN_828 : _GEN_827; // @[lut_mem_online.scala 234:34]
  wire  _GEN_830 = ~io_inputBit ? 1'h0 : _GEN_829; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_831 = i == 8'h50 ? _GEN_830 : _GEN_829; // @[lut_mem_online.scala 234:34]
  wire  _GEN_832 = io_inputBit | _GEN_831; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_833 = i == 8'h50 ? _GEN_832 : _GEN_831; // @[lut_mem_online.scala 234:34]
  wire  _GEN_834 = io_inputBit ? 1'h0 : _GEN_833; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_835 = i == 8'h51 ? _GEN_834 : _GEN_833; // @[lut_mem_online.scala 234:34]
  wire  _GEN_836 = io_inputBit | _GEN_835; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_837 = i == 8'h58 ? _GEN_836 : _GEN_835; // @[lut_mem_online.scala 234:34]
  wire  _GEN_838 = io_inputBit ? 1'h0 : _GEN_837; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_839 = i == 8'h59 ? _GEN_838 : _GEN_837; // @[lut_mem_online.scala 234:34]
  wire  _GEN_840 = ~io_inputBit | _GEN_839; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_841 = i == 8'h5a ? _GEN_840 : _GEN_839; // @[lut_mem_online.scala 234:34]
  wire  _GEN_842 = ~io_inputBit ? 1'h0 : _GEN_841; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_843 = i == 8'h5b ? _GEN_842 : _GEN_841; // @[lut_mem_online.scala 234:34]
  wire  _GEN_844 = io_inputBit | _GEN_843; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_845 = i == 8'h5b ? _GEN_844 : _GEN_843; // @[lut_mem_online.scala 234:34]
  wire  _GEN_846 = io_inputBit ? 1'h0 : _GEN_845; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_847 = i == 8'h5c ? _GEN_846 : _GEN_845; // @[lut_mem_online.scala 234:34]
  wire  _GEN_848 = ~io_inputBit | _GEN_847; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_849 = i == 8'ha0 ? _GEN_848 : _GEN_847; // @[lut_mem_online.scala 234:34]
  wire  _GEN_850 = io_inputBit ? 1'h0 : _GEN_849; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_851 = i == 8'ha0 ? _GEN_850 : _GEN_849; // @[lut_mem_online.scala 234:34]
  wire  _GEN_852 = ~io_inputBit | _GEN_851; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_853 = i == 8'ha3 ? _GEN_852 : _GEN_851; // @[lut_mem_online.scala 234:34]
  wire  _GEN_854 = io_inputBit ? 1'h0 : _GEN_853; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_855 = i == 8'ha3 ? _GEN_854 : _GEN_853; // @[lut_mem_online.scala 234:34]
  wire  _GEN_856 = ~io_inputBit ? 1'h0 : _GEN_855; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_857 = i == 8'hb1 ? _GEN_856 : _GEN_855; // @[lut_mem_online.scala 234:34]
  wire  _GEN_858 = io_inputBit | _GEN_857; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_859 = i == 8'hb1 ? _GEN_858 : _GEN_857; // @[lut_mem_online.scala 234:34]
  wire  _GEN_860 = ~io_inputBit | _GEN_859; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_861 = i == 8'hb3 ? _GEN_860 : _GEN_859; // @[lut_mem_online.scala 234:34]
  wire  _GEN_862 = io_inputBit ? 1'h0 : _GEN_861; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_863 = i == 8'hb3 ? _GEN_862 : _GEN_861; // @[lut_mem_online.scala 234:34]
  wire  _GEN_864 = ~io_inputBit | _GEN_863; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_865 = i == 8'hb6 ? _GEN_864 : _GEN_863; // @[lut_mem_online.scala 234:34]
  wire  _GEN_866 = io_inputBit ? 1'h0 : _GEN_865; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_867 = i == 8'hb6 ? _GEN_866 : _GEN_865; // @[lut_mem_online.scala 234:34]
  wire  _GEN_868 = ~io_inputBit | _GEN_867; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_869 = i == 8'hb9 ? _GEN_868 : _GEN_867; // @[lut_mem_online.scala 234:34]
  wire  _GEN_870 = io_inputBit ? 1'h0 : _GEN_869; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_871 = i == 8'hb9 ? _GEN_870 : _GEN_869; // @[lut_mem_online.scala 234:34]
  wire  _GEN_872 = io_inputBit ? 1'h0 : _GEN_491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_873 = i == 8'h0 ? _GEN_872 : _GEN_491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_874 = ~io_inputBit ? 1'h0 : _GEN_873; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_875 = i == 8'h3 ? _GEN_874 : _GEN_873; // @[lut_mem_online.scala 234:34]
  wire  _GEN_876 = ~io_inputBit ? 1'h0 : _GEN_875; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_877 = i == 8'h8 ? _GEN_876 : _GEN_875; // @[lut_mem_online.scala 234:34]
  wire  _GEN_878 = io_inputBit ? 1'h0 : _GEN_877; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_879 = i == 8'h9 ? _GEN_878 : _GEN_877; // @[lut_mem_online.scala 234:34]
  wire  _GEN_880 = ~io_inputBit ? 1'h0 : _GEN_879; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_881 = i == 8'h12 ? _GEN_880 : _GEN_879; // @[lut_mem_online.scala 234:34]
  wire  _GEN_882 = io_inputBit ? 1'h0 : _GEN_881; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_883 = i == 8'h16 ? _GEN_882 : _GEN_881; // @[lut_mem_online.scala 234:34]
  wire  _GEN_884 = ~io_inputBit ? 1'h0 : _GEN_883; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_885 = i == 8'h26 ? _GEN_884 : _GEN_883; // @[lut_mem_online.scala 234:34]
  wire  _GEN_886 = ~io_inputBit ? 1'h0 : _GEN_885; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_887 = i == 8'h2b ? _GEN_886 : _GEN_885; // @[lut_mem_online.scala 234:34]
  wire  _GEN_888 = ~io_inputBit ? 1'h0 : _GEN_887; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_889 = i == 8'h4e ? _GEN_888 : _GEN_887; // @[lut_mem_online.scala 234:34]
  wire  _GEN_890 = io_inputBit | _GEN_889; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_891 = i == 8'h4e ? _GEN_890 : _GEN_889; // @[lut_mem_online.scala 234:34]
  wire  _GEN_892 = ~io_inputBit | _GEN_891; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_893 = i == 8'h50 ? _GEN_892 : _GEN_891; // @[lut_mem_online.scala 234:34]
  wire  _GEN_894 = io_inputBit ? 1'h0 : _GEN_893; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_895 = i == 8'h50 ? _GEN_894 : _GEN_893; // @[lut_mem_online.scala 234:34]
  wire  _GEN_896 = ~io_inputBit ? 1'h0 : _GEN_895; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_897 = i == 8'h52 ? _GEN_896 : _GEN_895; // @[lut_mem_online.scala 234:34]
  wire  _GEN_898 = io_inputBit | _GEN_897; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_899 = i == 8'h52 ? _GEN_898 : _GEN_897; // @[lut_mem_online.scala 234:34]
  wire  _GEN_900 = io_inputBit ? 1'h0 : _GEN_899; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_901 = i == 8'h59 ? _GEN_900 : _GEN_899; // @[lut_mem_online.scala 234:34]
  wire  _GEN_902 = io_inputBit | _GEN_901; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_903 = i == 8'h5b ? _GEN_902 : _GEN_901; // @[lut_mem_online.scala 234:34]
  wire  _GEN_904 = ~io_inputBit ? 1'h0 : _GEN_903; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_905 = i == 8'h9f ? _GEN_904 : _GEN_903; // @[lut_mem_online.scala 234:34]
  wire  _GEN_906 = io_inputBit | _GEN_905; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_907 = i == 8'h9f ? _GEN_906 : _GEN_905; // @[lut_mem_online.scala 234:34]
  wire  _GEN_908 = ~io_inputBit | _GEN_907; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_909 = i == 8'ha0 ? _GEN_908 : _GEN_907; // @[lut_mem_online.scala 234:34]
  wire  _GEN_910 = io_inputBit ? 1'h0 : _GEN_909; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_911 = i == 8'ha0 ? _GEN_910 : _GEN_909; // @[lut_mem_online.scala 234:34]
  wire  _GEN_912 = ~io_inputBit | _GEN_911; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_913 = i == 8'ha3 ? _GEN_912 : _GEN_911; // @[lut_mem_online.scala 234:34]
  wire  _GEN_914 = io_inputBit ? 1'h0 : _GEN_913; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_915 = i == 8'ha3 ? _GEN_914 : _GEN_913; // @[lut_mem_online.scala 234:34]
  wire  _GEN_916 = ~io_inputBit ? 1'h0 : _GEN_915; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_917 = i == 8'ha4 ? _GEN_916 : _GEN_915; // @[lut_mem_online.scala 234:34]
  wire  _GEN_918 = io_inputBit | _GEN_917; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_919 = i == 8'ha4 ? _GEN_918 : _GEN_917; // @[lut_mem_online.scala 234:34]
  wire  _GEN_920 = ~io_inputBit ? 1'h0 : _GEN_919; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_921 = i == 8'hb1 ? _GEN_920 : _GEN_919; // @[lut_mem_online.scala 234:34]
  wire  _GEN_922 = io_inputBit | _GEN_921; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_923 = i == 8'hb1 ? _GEN_922 : _GEN_921; // @[lut_mem_online.scala 234:34]
  wire  _GEN_924 = ~io_inputBit | _GEN_923; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_925 = i == 8'hb2 ? _GEN_924 : _GEN_923; // @[lut_mem_online.scala 234:34]
  wire  _GEN_926 = io_inputBit ? 1'h0 : _GEN_925; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_927 = i == 8'hb2 ? _GEN_926 : _GEN_925; // @[lut_mem_online.scala 234:34]
  wire  _GEN_928 = ~io_inputBit ? 1'h0 : _GEN_927; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_929 = i == 8'hb3 ? _GEN_928 : _GEN_927; // @[lut_mem_online.scala 234:34]
  wire  _GEN_930 = io_inputBit | _GEN_929; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_931 = i == 8'hb3 ? _GEN_930 : _GEN_929; // @[lut_mem_online.scala 234:34]
  wire  _GEN_932 = ~io_inputBit | _GEN_931; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_933 = i == 8'hb5 ? _GEN_932 : _GEN_931; // @[lut_mem_online.scala 234:34]
  wire  _GEN_934 = io_inputBit ? 1'h0 : _GEN_933; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_935 = i == 8'hb5 ? _GEN_934 : _GEN_933; // @[lut_mem_online.scala 234:34]
  wire  _GEN_936 = ~io_inputBit ? 1'h0 : _GEN_935; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_937 = i == 8'hb6 ? _GEN_936 : _GEN_935; // @[lut_mem_online.scala 234:34]
  wire  _GEN_938 = io_inputBit | _GEN_937; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_939 = i == 8'hb6 ? _GEN_938 : _GEN_937; // @[lut_mem_online.scala 234:34]
  wire  _GEN_940 = ~io_inputBit | _GEN_939; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_941 = i == 8'hb7 ? _GEN_940 : _GEN_939; // @[lut_mem_online.scala 234:34]
  wire  _GEN_942 = io_inputBit ? 1'h0 : _GEN_941; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_943 = i == 8'hb7 ? _GEN_942 : _GEN_941; // @[lut_mem_online.scala 234:34]
  wire  _GEN_944 = ~io_inputBit ? 1'h0 : _GEN_943; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_945 = i == 8'hb9 ? _GEN_944 : _GEN_943; // @[lut_mem_online.scala 234:34]
  wire  _GEN_946 = io_inputBit | _GEN_945; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_947 = i == 8'hb9 ? _GEN_946 : _GEN_945; // @[lut_mem_online.scala 234:34]
  wire  _GEN_948 = ~io_inputBit | _GEN_947; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_949 = i == 8'hba ? _GEN_948 : _GEN_947; // @[lut_mem_online.scala 234:34]
  wire  _GEN_950 = io_inputBit ? 1'h0 : _GEN_949; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_951 = i == 8'hba ? _GEN_950 : _GEN_949; // @[lut_mem_online.scala 234:34]
  wire  _GEN_952 = io_inputBit ? 1'h0 : _GEN_577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_953 = i == 8'h0 ? _GEN_952 : _GEN_577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_954 = ~io_inputBit ? 1'h0 : _GEN_953; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_955 = i == 8'h3 ? _GEN_954 : _GEN_953; // @[lut_mem_online.scala 234:34]
  wire  _GEN_956 = ~io_inputBit ? 1'h0 : _GEN_955; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_957 = i == 8'h8 ? _GEN_956 : _GEN_955; // @[lut_mem_online.scala 234:34]
  wire  _GEN_958 = io_inputBit | _GEN_957; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_959 = i == 8'h9 ? _GEN_958 : _GEN_957; // @[lut_mem_online.scala 234:34]
  wire  _GEN_960 = ~io_inputBit ? 1'h0 : _GEN_959; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_961 = i == 8'h12 ? _GEN_960 : _GEN_959; // @[lut_mem_online.scala 234:34]
  wire  _GEN_962 = io_inputBit ? 1'h0 : _GEN_961; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_963 = i == 8'h16 ? _GEN_962 : _GEN_961; // @[lut_mem_online.scala 234:34]
  wire  _GEN_964 = ~io_inputBit ? 1'h0 : _GEN_963; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_965 = i == 8'h26 ? _GEN_964 : _GEN_963; // @[lut_mem_online.scala 234:34]
  wire  _GEN_966 = ~io_inputBit | _GEN_965; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_967 = i == 8'h2b ? _GEN_966 : _GEN_965; // @[lut_mem_online.scala 234:34]
  wire  _GEN_968 = ~io_inputBit | _GEN_967; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_969 = i == 8'h58 ? _GEN_968 : _GEN_967; // @[lut_mem_online.scala 234:34]
  wire  _GEN_970 = ~io_inputBit ? 1'h0 : _GEN_969; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_971 = i == 8'h59 ? _GEN_970 : _GEN_969; // @[lut_mem_online.scala 234:34]
  wire  _GEN_972 = ~io_inputBit | _GEN_971; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_973 = i == 8'h5a ? _GEN_972 : _GEN_971; // @[lut_mem_online.scala 234:34]
  wire  _GEN_974 = ~io_inputBit ? 1'h0 : _GEN_973; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_975 = i == 8'h5b ? _GEN_974 : _GEN_973; // @[lut_mem_online.scala 234:34]
  wire  _GEN_976 = ~io_inputBit | _GEN_975; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_977 = i == 8'h5c ? _GEN_976 : _GEN_975; // @[lut_mem_online.scala 234:34]
  wire  _GEN_978 = ~io_inputBit ? 1'h0 : _GEN_977; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_979 = i == 8'h9d ? _GEN_978 : _GEN_977; // @[lut_mem_online.scala 234:34]
  wire  _GEN_980 = io_inputBit | _GEN_979; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_981 = i == 8'h9d ? _GEN_980 : _GEN_979; // @[lut_mem_online.scala 234:34]
  wire  _GEN_982 = ~io_inputBit ? 1'h0 : _GEN_981; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_983 = i == 8'h9e ? _GEN_982 : _GEN_981; // @[lut_mem_online.scala 234:34]
  wire  _GEN_984 = io_inputBit | _GEN_983; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_985 = i == 8'h9e ? _GEN_984 : _GEN_983; // @[lut_mem_online.scala 234:34]
  wire  _GEN_986 = ~io_inputBit | _GEN_985; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_987 = i == 8'h9f ? _GEN_986 : _GEN_985; // @[lut_mem_online.scala 234:34]
  wire  _GEN_988 = io_inputBit ? 1'h0 : _GEN_987; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_989 = i == 8'h9f ? _GEN_988 : _GEN_987; // @[lut_mem_online.scala 234:34]
  wire  _GEN_990 = ~io_inputBit | _GEN_989; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_991 = i == 8'ha0 ? _GEN_990 : _GEN_989; // @[lut_mem_online.scala 234:34]
  wire  _GEN_992 = io_inputBit ? 1'h0 : _GEN_991; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_993 = i == 8'ha0 ? _GEN_992 : _GEN_991; // @[lut_mem_online.scala 234:34]
  wire  _GEN_994 = ~io_inputBit ? 1'h0 : _GEN_993; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_995 = i == 8'ha1 ? _GEN_994 : _GEN_993; // @[lut_mem_online.scala 234:34]
  wire  _GEN_996 = io_inputBit | _GEN_995; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_997 = i == 8'ha1 ? _GEN_996 : _GEN_995; // @[lut_mem_online.scala 234:34]
  wire  _GEN_998 = ~io_inputBit ? 1'h0 : _GEN_997; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_999 = i == 8'ha2 ? _GEN_998 : _GEN_997; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1000 = io_inputBit | _GEN_999; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1001 = i == 8'ha2 ? _GEN_1000 : _GEN_999; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1002 = ~io_inputBit | _GEN_1001; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1003 = i == 8'ha3 ? _GEN_1002 : _GEN_1001; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1004 = io_inputBit ? 1'h0 : _GEN_1003; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1005 = i == 8'ha3 ? _GEN_1004 : _GEN_1003; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1006 = ~io_inputBit | _GEN_1005; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1007 = i == 8'ha4 ? _GEN_1006 : _GEN_1005; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1008 = io_inputBit ? 1'h0 : _GEN_1007; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1009 = i == 8'ha4 ? _GEN_1008 : _GEN_1007; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1010 = ~io_inputBit ? 1'h0 : _GEN_1009; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1011 = i == 8'ha5 ? _GEN_1010 : _GEN_1009; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1012 = io_inputBit | _GEN_1011; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1013 = i == 8'ha5 ? _GEN_1012 : _GEN_1011; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1014 = ~io_inputBit ? 1'h0 : _GEN_1013; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1015 = i == 8'ha6 ? _GEN_1014 : _GEN_1013; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1016 = io_inputBit | _GEN_1015; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1017 = i == 8'ha6 ? _GEN_1016 : _GEN_1015; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1018 = ~io_inputBit ? 1'h0 : _GEN_1017; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1019 = i == 8'hb2 ? _GEN_1018 : _GEN_1017; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1020 = io_inputBit | _GEN_1019; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1021 = i == 8'hb2 ? _GEN_1020 : _GEN_1019; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1022 = ~io_inputBit | _GEN_1021; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1023 = i == 8'hb4 ? _GEN_1022 : _GEN_1021; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1024 = io_inputBit ? 1'h0 : _GEN_1023; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1025 = i == 8'hb4 ? _GEN_1024 : _GEN_1023; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1026 = ~io_inputBit ? 1'h0 : _GEN_1025; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1027 = i == 8'hb6 ? _GEN_1026 : _GEN_1025; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1028 = io_inputBit | _GEN_1027; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1029 = i == 8'hb6 ? _GEN_1028 : _GEN_1027; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1030 = ~io_inputBit | _GEN_1029; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1031 = i == 8'hb8 ? _GEN_1030 : _GEN_1029; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1032 = io_inputBit ? 1'h0 : _GEN_1031; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1033 = i == 8'hb8 ? _GEN_1032 : _GEN_1031; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1034 = ~io_inputBit ? 1'h0 : _GEN_1033; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1035 = i == 8'hba ? _GEN_1034 : _GEN_1033; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1036 = io_inputBit | _GEN_1035; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1037 = i == 8'hba ? _GEN_1036 : _GEN_1035; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1038 = io_inputBit ? 1'h0 : _GEN_653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1039 = i == 8'h0 ? _GEN_1038 : _GEN_653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1040 = ~io_inputBit ? 1'h0 : _GEN_1039; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1041 = i == 8'h3 ? _GEN_1040 : _GEN_1039; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1042 = ~io_inputBit ? 1'h0 : _GEN_1041; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1043 = i == 8'h8 ? _GEN_1042 : _GEN_1041; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1044 = io_inputBit ? 1'h0 : _GEN_1043; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1045 = i == 8'h9 ? _GEN_1044 : _GEN_1043; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1046 = ~io_inputBit ? 1'h0 : _GEN_1045; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1047 = i == 8'h12 ? _GEN_1046 : _GEN_1045; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1048 = io_inputBit ? 1'h0 : _GEN_1047; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1049 = i == 8'h16 ? _GEN_1048 : _GEN_1047; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1050 = ~io_inputBit ? 1'h0 : _GEN_1049; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1051 = i == 8'h26 ? _GEN_1050 : _GEN_1049; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1052 = ~io_inputBit ? 1'h0 : _GEN_1051; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1053 = i == 8'h2b ? _GEN_1052 : _GEN_1051; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1054 = ~io_inputBit ? 1'h0 : _GEN_1053; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1055 = i == 8'h4e ? _GEN_1054 : _GEN_1053; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1056 = io_inputBit | _GEN_1055; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1057 = i == 8'h4e ? _GEN_1056 : _GEN_1055; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1058 = ~io_inputBit ? 1'h0 : _GEN_1057; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1059 = i == 8'h4f ? _GEN_1058 : _GEN_1057; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1060 = io_inputBit | _GEN_1059; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1061 = i == 8'h4f ? _GEN_1060 : _GEN_1059; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1062 = ~io_inputBit ? 1'h0 : _GEN_1061; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1063 = i == 8'h50 ? _GEN_1062 : _GEN_1061; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1064 = io_inputBit | _GEN_1063; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1065 = i == 8'h50 ? _GEN_1064 : _GEN_1063; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1066 = ~io_inputBit ? 1'h0 : _GEN_1065; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1067 = i == 8'h51 ? _GEN_1066 : _GEN_1065; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1068 = io_inputBit | _GEN_1067; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1069 = i == 8'h51 ? _GEN_1068 : _GEN_1067; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1070 = ~io_inputBit ? 1'h0 : _GEN_1069; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1071 = i == 8'h52 ? _GEN_1070 : _GEN_1069; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1072 = io_inputBit | _GEN_1071; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1073 = i == 8'h52 ? _GEN_1072 : _GEN_1071; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1074 = ~io_inputBit ? 1'h0 : _GEN_1073; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1075 = i == 8'hb1 ? _GEN_1074 : _GEN_1073; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1076 = io_inputBit | _GEN_1075; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1077 = i == 8'hb1 ? _GEN_1076 : _GEN_1075; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1078 = ~io_inputBit | _GEN_1077; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1079 = i == 8'hb2 ? _GEN_1078 : _GEN_1077; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1080 = io_inputBit ? 1'h0 : _GEN_1079; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1081 = i == 8'hb2 ? _GEN_1080 : _GEN_1079; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1082 = ~io_inputBit ? 1'h0 : _GEN_1081; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1083 = i == 8'hb3 ? _GEN_1082 : _GEN_1081; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1084 = io_inputBit | _GEN_1083; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1085 = i == 8'hb3 ? _GEN_1084 : _GEN_1083; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1086 = ~io_inputBit | _GEN_1085; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1087 = i == 8'hb4 ? _GEN_1086 : _GEN_1085; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1088 = io_inputBit ? 1'h0 : _GEN_1087; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1089 = i == 8'hb4 ? _GEN_1088 : _GEN_1087; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1090 = ~io_inputBit ? 1'h0 : _GEN_1089; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1091 = i == 8'hb5 ? _GEN_1090 : _GEN_1089; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1092 = io_inputBit | _GEN_1091; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1093 = i == 8'hb5 ? _GEN_1092 : _GEN_1091; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1094 = ~io_inputBit | _GEN_1093; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1095 = i == 8'hb6 ? _GEN_1094 : _GEN_1093; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1096 = io_inputBit ? 1'h0 : _GEN_1095; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1097 = i == 8'hb6 ? _GEN_1096 : _GEN_1095; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1098 = ~io_inputBit ? 1'h0 : _GEN_1097; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1099 = i == 8'hb7 ? _GEN_1098 : _GEN_1097; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1100 = io_inputBit | _GEN_1099; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1101 = i == 8'hb7 ? _GEN_1100 : _GEN_1099; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1102 = ~io_inputBit | _GEN_1101; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1103 = i == 8'hb8 ? _GEN_1102 : _GEN_1101; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1104 = io_inputBit ? 1'h0 : _GEN_1103; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1105 = i == 8'hb8 ? _GEN_1104 : _GEN_1103; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1106 = ~io_inputBit ? 1'h0 : _GEN_1105; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1107 = i == 8'hb9 ? _GEN_1106 : _GEN_1105; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1108 = io_inputBit | _GEN_1107; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1109 = i == 8'hb9 ? _GEN_1108 : _GEN_1107; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1110 = ~io_inputBit | _GEN_1109; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1111 = i == 8'hba ? _GEN_1110 : _GEN_1109; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1112 = io_inputBit ? 1'h0 : _GEN_1111; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1113 = i == 8'hba ? _GEN_1112 : _GEN_1111; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1114 = io_inputBit ? 1'h0 : _GEN_749; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1115 = i == 8'h0 ? _GEN_1114 : _GEN_749; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1116 = ~io_inputBit ? 1'h0 : _GEN_1115; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1117 = i == 8'h3 ? _GEN_1116 : _GEN_1115; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1118 = ~io_inputBit ? 1'h0 : _GEN_1117; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1119 = i == 8'h8 ? _GEN_1118 : _GEN_1117; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1120 = io_inputBit ? 1'h0 : _GEN_1119; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1121 = i == 8'h9 ? _GEN_1120 : _GEN_1119; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1122 = ~io_inputBit ? 1'h0 : _GEN_1121; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1123 = i == 8'h12 ? _GEN_1122 : _GEN_1121; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1124 = io_inputBit ? 1'h0 : _GEN_1123; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1125 = i == 8'h16 ? _GEN_1124 : _GEN_1123; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1126 = ~io_inputBit ? 1'h0 : _GEN_1125; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1127 = i == 8'h26 ? _GEN_1126 : _GEN_1125; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1128 = ~io_inputBit ? 1'h0 : _GEN_1127; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1129 = i == 8'h2b ? _GEN_1128 : _GEN_1127; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1130 = ~io_inputBit ? 1'h0 : _GEN_1129; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1131 = i == 8'h9d ? _GEN_1130 : _GEN_1129; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1132 = io_inputBit | _GEN_1131; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1133 = i == 8'h9d ? _GEN_1132 : _GEN_1131; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1134 = ~io_inputBit ? 1'h0 : _GEN_1133; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1135 = i == 8'h9e ? _GEN_1134 : _GEN_1133; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1136 = io_inputBit | _GEN_1135; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1137 = i == 8'h9e ? _GEN_1136 : _GEN_1135; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1138 = ~io_inputBit ? 1'h0 : _GEN_1137; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1139 = i == 8'h9f ? _GEN_1138 : _GEN_1137; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1140 = io_inputBit | _GEN_1139; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1141 = i == 8'h9f ? _GEN_1140 : _GEN_1139; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1142 = ~io_inputBit ? 1'h0 : _GEN_1141; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1143 = i == 8'ha0 ? _GEN_1142 : _GEN_1141; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1144 = io_inputBit | _GEN_1143; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1145 = i == 8'ha0 ? _GEN_1144 : _GEN_1143; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1146 = ~io_inputBit ? 1'h0 : _GEN_1145; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1147 = i == 8'ha1 ? _GEN_1146 : _GEN_1145; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1148 = io_inputBit | _GEN_1147; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1149 = i == 8'ha1 ? _GEN_1148 : _GEN_1147; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1150 = ~io_inputBit ? 1'h0 : _GEN_1149; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1151 = i == 8'ha2 ? _GEN_1150 : _GEN_1149; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1152 = io_inputBit | _GEN_1151; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1153 = i == 8'ha2 ? _GEN_1152 : _GEN_1151; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1154 = ~io_inputBit ? 1'h0 : _GEN_1153; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1155 = i == 8'ha3 ? _GEN_1154 : _GEN_1153; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1156 = io_inputBit | _GEN_1155; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1157 = i == 8'ha3 ? _GEN_1156 : _GEN_1155; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1158 = ~io_inputBit ? 1'h0 : _GEN_1157; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1159 = i == 8'ha4 ? _GEN_1158 : _GEN_1157; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1160 = io_inputBit | _GEN_1159; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1161 = i == 8'ha4 ? _GEN_1160 : _GEN_1159; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1162 = ~io_inputBit ? 1'h0 : _GEN_1161; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1163 = i == 8'ha5 ? _GEN_1162 : _GEN_1161; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1164 = io_inputBit | _GEN_1163; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1165 = i == 8'ha5 ? _GEN_1164 : _GEN_1163; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1166 = ~io_inputBit ? 1'h0 : _GEN_1165; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1167 = i == 8'ha6 ? _GEN_1166 : _GEN_1165; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1168 = io_inputBit | _GEN_1167; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1169 = i == 8'ha6 ? _GEN_1168 : _GEN_1167; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1170 = ~io_inputBit ? 1'h0 : _GEN_1169; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1171 = i == 8'hb1 ? _GEN_1170 : _GEN_1169; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1172 = io_inputBit | _GEN_1171; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1173 = i == 8'hb1 ? _GEN_1172 : _GEN_1171; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1174 = ~io_inputBit ? 1'h0 : _GEN_1173; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1175 = i == 8'hb2 ? _GEN_1174 : _GEN_1173; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1176 = io_inputBit | _GEN_1175; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1177 = i == 8'hb2 ? _GEN_1176 : _GEN_1175; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1178 = ~io_inputBit ? 1'h0 : _GEN_1177; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1179 = i == 8'hb3 ? _GEN_1178 : _GEN_1177; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1180 = io_inputBit | _GEN_1179; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1181 = i == 8'hb3 ? _GEN_1180 : _GEN_1179; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1182 = ~io_inputBit ? 1'h0 : _GEN_1181; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1183 = i == 8'hb4 ? _GEN_1182 : _GEN_1181; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1184 = io_inputBit | _GEN_1183; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1185 = i == 8'hb4 ? _GEN_1184 : _GEN_1183; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1186 = ~io_inputBit ? 1'h0 : _GEN_1185; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1187 = i == 8'hb5 ? _GEN_1186 : _GEN_1185; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1188 = io_inputBit | _GEN_1187; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1189 = i == 8'hb5 ? _GEN_1188 : _GEN_1187; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1190 = ~io_inputBit ? 1'h0 : _GEN_1189; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1191 = i == 8'hb6 ? _GEN_1190 : _GEN_1189; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1192 = io_inputBit | _GEN_1191; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1193 = i == 8'hb6 ? _GEN_1192 : _GEN_1191; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1194 = ~io_inputBit ? 1'h0 : _GEN_1193; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1195 = i == 8'hb7 ? _GEN_1194 : _GEN_1193; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1196 = io_inputBit | _GEN_1195; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1197 = i == 8'hb7 ? _GEN_1196 : _GEN_1195; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1198 = ~io_inputBit ? 1'h0 : _GEN_1197; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1199 = i == 8'hb8 ? _GEN_1198 : _GEN_1197; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1200 = io_inputBit | _GEN_1199; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1201 = i == 8'hb8 ? _GEN_1200 : _GEN_1199; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1202 = ~io_inputBit ? 1'h0 : _GEN_1201; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1203 = i == 8'hb9 ? _GEN_1202 : _GEN_1201; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1204 = io_inputBit | _GEN_1203; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1205 = i == 8'hb9 ? _GEN_1204 : _GEN_1203; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1206 = ~io_inputBit ? 1'h0 : _GEN_1205; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1207 = i == 8'hba ? _GEN_1206 : _GEN_1205; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1208 = io_inputBit | _GEN_1207; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1209 = i == 8'hba ? _GEN_1208 : _GEN_1207; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1210 = ~io_inputBit ? 1'h0 : _GEN_773; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1211 = i == 8'h1 ? _GEN_1210 : _GEN_773; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1212 = io_inputBit ? 1'h0 : _GEN_1211; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1213 = i == 8'h2 ? _GEN_1212 : _GEN_1211; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1214 = ~io_inputBit ? 1'h0 : _GEN_1213; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1215 = i == 8'h4 ? _GEN_1214 : _GEN_1213; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1216 = io_inputBit ? 1'h0 : _GEN_1215; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1217 = i == 8'h5 ? _GEN_1216 : _GEN_1215; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1218 = ~io_inputBit ? 1'h0 : _GEN_1217; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1219 = i == 8'ha ? _GEN_1218 : _GEN_1217; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1220 = ~io_inputBit | _GEN_1219; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1221 = i == 8'hb ? _GEN_1220 : _GEN_1219; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1222 = io_inputBit | _GEN_1221; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1223 = i == 8'h16 ? _GEN_1222 : _GEN_1221; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1224 = io_inputBit ? 1'h0 : _GEN_1223; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1225 = i == 8'h18 ? _GEN_1224 : _GEN_1223; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1226 = io_inputBit | _GEN_1225; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1227 = i == 8'h2d ? _GEN_1226 : _GEN_1225; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1228 = ~io_inputBit | _GEN_1227; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1229 = i == 8'h31 ? _GEN_1228 : _GEN_1227; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1230 = io_inputBit ? 1'h0 : _GEN_1229; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1231 = i == 8'h31 ? _GEN_1230 : _GEN_1229; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1232 = io_inputBit | _GEN_1231; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1233 = i == 8'h5b ? _GEN_1232 : _GEN_1231; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1234 = ~io_inputBit ? 1'h0 : _GEN_1233; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1235 = i == 8'hb7 ? _GEN_1234 : _GEN_1233; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1236 = io_inputBit | _GEN_1235; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1238 = ~io_inputBit ? 1'h0 : _GEN_815; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1239 = i == 8'h1 ? _GEN_1238 : _GEN_815; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1240 = io_inputBit ? 1'h0 : _GEN_1239; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1241 = i == 8'h2 ? _GEN_1240 : _GEN_1239; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1242 = ~io_inputBit ? 1'h0 : _GEN_1241; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1243 = i == 8'h4 ? _GEN_1242 : _GEN_1241; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1244 = io_inputBit ? 1'h0 : _GEN_1243; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1245 = i == 8'h5 ? _GEN_1244 : _GEN_1243; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1246 = ~io_inputBit ? 1'h0 : _GEN_1245; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1247 = i == 8'h15 ? _GEN_1246 : _GEN_1245; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1248 = io_inputBit | _GEN_1247; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1249 = i == 8'h16 ? _GEN_1248 : _GEN_1247; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1250 = ~io_inputBit | _GEN_1249; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1251 = i == 8'h17 ? _GEN_1250 : _GEN_1249; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1252 = io_inputBit | _GEN_1251; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1253 = i == 8'h2c ? _GEN_1252 : _GEN_1251; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1254 = io_inputBit ? 1'h0 : _GEN_1253; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1255 = i == 8'h2d ? _GEN_1254 : _GEN_1253; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1256 = ~io_inputBit | _GEN_1255; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1257 = i == 8'h30 ? _GEN_1256 : _GEN_1255; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1258 = ~io_inputBit ? 1'h0 : _GEN_1257; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1259 = i == 8'h31 ? _GEN_1258 : _GEN_1257; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1260 = io_inputBit | _GEN_1259; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1261 = i == 8'h31 ? _GEN_1260 : _GEN_1259; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1262 = io_inputBit ? 1'h0 : _GEN_1261; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1263 = i == 8'h32 ? _GEN_1262 : _GEN_1261; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1264 = ~io_inputBit ? 1'h0 : _GEN_1263; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1265 = i == 8'h59 ? _GEN_1264 : _GEN_1263; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1266 = io_inputBit ? 1'h0 : _GEN_1265; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1267 = i == 8'h5b ? _GEN_1266 : _GEN_1265; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1268 = io_inputBit ? 1'h0 : _GEN_1267; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1269 = i == 8'h62 ? _GEN_1268 : _GEN_1267; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1270 = ~io_inputBit | _GEN_1269; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1271 = i == 8'h65 ? _GEN_1270 : _GEN_1269; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1272 = io_inputBit ? 1'h0 : _GEN_1271; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1273 = i == 8'h65 ? _GEN_1272 : _GEN_1271; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1274 = ~io_inputBit ? 1'h0 : _GEN_1273; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1275 = i == 8'hb4 ? _GEN_1274 : _GEN_1273; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1276 = io_inputBit | _GEN_1275; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1277 = i == 8'hb4 ? _GEN_1276 : _GEN_1275; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1278 = ~io_inputBit | _GEN_1277; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1279 = i == 8'hb7 ? _GEN_1278 : _GEN_1277; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1280 = io_inputBit ? 1'h0 : _GEN_1279; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1281 = i == 8'hb7 ? _GEN_1280 : _GEN_1279; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1282 = ~io_inputBit | _GEN_1281; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1283 = i == 8'hc5 ? _GEN_1282 : _GEN_1281; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1286 = ~io_inputBit ? 1'h0 : _GEN_871; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1287 = i == 8'h1 ? _GEN_1286 : _GEN_871; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1288 = io_inputBit ? 1'h0 : _GEN_1287; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1289 = i == 8'h2 ? _GEN_1288 : _GEN_1287; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1290 = ~io_inputBit ? 1'h0 : _GEN_1289; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1291 = i == 8'h4 ? _GEN_1290 : _GEN_1289; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1292 = io_inputBit ? 1'h0 : _GEN_1291; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1293 = i == 8'h5 ? _GEN_1292 : _GEN_1291; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1294 = ~io_inputBit ? 1'h0 : _GEN_1293; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1295 = i == 8'h15 ? _GEN_1294 : _GEN_1293; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1296 = io_inputBit ? 1'h0 : _GEN_1295; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1297 = i == 8'h16 ? _GEN_1296 : _GEN_1295; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1298 = ~io_inputBit ? 1'h0 : _GEN_1297; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1299 = i == 8'h17 ? _GEN_1298 : _GEN_1297; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1300 = io_inputBit | _GEN_1299; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1301 = i == 8'h2d ? _GEN_1300 : _GEN_1299; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1302 = ~io_inputBit ? 1'h0 : _GEN_1301; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1303 = i == 8'h30 ? _GEN_1302 : _GEN_1301; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1304 = ~io_inputBit | _GEN_1303; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1305 = i == 8'h59 ? _GEN_1304 : _GEN_1303; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1306 = ~io_inputBit ? 1'h0 : _GEN_1305; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1307 = i == 8'h5a ? _GEN_1306 : _GEN_1305; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1308 = io_inputBit | _GEN_1307; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1309 = i == 8'h5a ? _GEN_1308 : _GEN_1307; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1310 = io_inputBit ? 1'h0 : _GEN_1309; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1311 = i == 8'h5b ? _GEN_1310 : _GEN_1309; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1312 = io_inputBit | _GEN_1311; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1313 = i == 8'h62 ? _GEN_1312 : _GEN_1311; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1314 = io_inputBit ? 1'h0 : _GEN_1313; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1315 = i == 8'h63 ? _GEN_1314 : _GEN_1313; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1316 = ~io_inputBit | _GEN_1315; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1317 = i == 8'h64 ? _GEN_1316 : _GEN_1315; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1318 = ~io_inputBit ? 1'h0 : _GEN_1317; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1319 = i == 8'h65 ? _GEN_1318 : _GEN_1317; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1320 = io_inputBit | _GEN_1319; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1321 = i == 8'h65 ? _GEN_1320 : _GEN_1319; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1322 = io_inputBit ? 1'h0 : _GEN_1321; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1323 = i == 8'h66 ? _GEN_1322 : _GEN_1321; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1324 = ~io_inputBit | _GEN_1323; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1325 = i == 8'hb4 ? _GEN_1324 : _GEN_1323; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1326 = io_inputBit ? 1'h0 : _GEN_1325; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1327 = i == 8'hb4 ? _GEN_1326 : _GEN_1325; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1328 = ~io_inputBit | _GEN_1327; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1329 = i == 8'hb7 ? _GEN_1328 : _GEN_1327; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1330 = io_inputBit ? 1'h0 : _GEN_1329; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1331 = i == 8'hb7 ? _GEN_1330 : _GEN_1329; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1332 = ~io_inputBit ? 1'h0 : _GEN_1331; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1333 = i == 8'hc5 ? _GEN_1332 : _GEN_1331; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1334 = io_inputBit | _GEN_1333; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1335 = i == 8'hc5 ? _GEN_1334 : _GEN_1333; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1336 = ~io_inputBit | _GEN_1335; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1337 = i == 8'hc7 ? _GEN_1336 : _GEN_1335; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1338 = io_inputBit ? 1'h0 : _GEN_1337; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1339 = i == 8'hc7 ? _GEN_1338 : _GEN_1337; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1340 = ~io_inputBit | _GEN_1339; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1341 = i == 8'hca ? _GEN_1340 : _GEN_1339; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1342 = io_inputBit ? 1'h0 : _GEN_1341; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1343 = i == 8'hca ? _GEN_1342 : _GEN_1341; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1344 = ~io_inputBit | _GEN_1343; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1345 = i == 8'hcd ? _GEN_1344 : _GEN_1343; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1348 = ~io_inputBit ? 1'h0 : _GEN_951; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1349 = i == 8'h1 ? _GEN_1348 : _GEN_951; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1350 = io_inputBit ? 1'h0 : _GEN_1349; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1351 = i == 8'h2 ? _GEN_1350 : _GEN_1349; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1352 = ~io_inputBit ? 1'h0 : _GEN_1351; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1353 = i == 8'h4 ? _GEN_1352 : _GEN_1351; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1354 = io_inputBit ? 1'h0 : _GEN_1353; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1355 = i == 8'h5 ? _GEN_1354 : _GEN_1353; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1356 = io_inputBit ? 1'h0 : _GEN_1355; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1357 = i == 8'h16 ? _GEN_1356 : _GEN_1355; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1358 = ~io_inputBit ? 1'h0 : _GEN_1357; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1359 = i == 8'h17 ? _GEN_1358 : _GEN_1357; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1360 = ~io_inputBit ? 1'h0 : _GEN_1359; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1361 = i == 8'h2b ? _GEN_1360 : _GEN_1359; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1362 = ~io_inputBit ? 1'h0 : _GEN_1361; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1363 = i == 8'h30 ? _GEN_1362 : _GEN_1361; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1364 = ~io_inputBit ? 1'h0 : _GEN_1363; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1365 = i == 8'h58 ? _GEN_1364 : _GEN_1363; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1366 = io_inputBit | _GEN_1365; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1367 = i == 8'h58 ? _GEN_1366 : _GEN_1365; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1368 = ~io_inputBit | _GEN_1367; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1369 = i == 8'h5a ? _GEN_1368 : _GEN_1367; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1370 = io_inputBit ? 1'h0 : _GEN_1369; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1371 = i == 8'h5a ? _GEN_1370 : _GEN_1369; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1372 = ~io_inputBit ? 1'h0 : _GEN_1371; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1373 = i == 8'h5c ? _GEN_1372 : _GEN_1371; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1374 = io_inputBit | _GEN_1373; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1375 = i == 8'h5c ? _GEN_1374 : _GEN_1373; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1376 = io_inputBit ? 1'h0 : _GEN_1375; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1377 = i == 8'h63 ? _GEN_1376 : _GEN_1375; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1378 = io_inputBit | _GEN_1377; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1379 = i == 8'h65 ? _GEN_1378 : _GEN_1377; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1380 = ~io_inputBit ? 1'h0 : _GEN_1379; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1381 = i == 8'hb3 ? _GEN_1380 : _GEN_1379; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1382 = io_inputBit | _GEN_1381; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1383 = i == 8'hb3 ? _GEN_1382 : _GEN_1381; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1384 = ~io_inputBit | _GEN_1383; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1385 = i == 8'hb4 ? _GEN_1384 : _GEN_1383; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1386 = io_inputBit ? 1'h0 : _GEN_1385; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1387 = i == 8'hb4 ? _GEN_1386 : _GEN_1385; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1388 = ~io_inputBit | _GEN_1387; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1389 = i == 8'hb7 ? _GEN_1388 : _GEN_1387; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1390 = io_inputBit ? 1'h0 : _GEN_1389; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1391 = i == 8'hb7 ? _GEN_1390 : _GEN_1389; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1392 = ~io_inputBit ? 1'h0 : _GEN_1391; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1393 = i == 8'hb8 ? _GEN_1392 : _GEN_1391; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1394 = io_inputBit | _GEN_1393; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1395 = i == 8'hb8 ? _GEN_1394 : _GEN_1393; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1396 = ~io_inputBit ? 1'h0 : _GEN_1395; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1397 = i == 8'hc5 ? _GEN_1396 : _GEN_1395; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1398 = io_inputBit | _GEN_1397; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1399 = i == 8'hc5 ? _GEN_1398 : _GEN_1397; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1400 = ~io_inputBit | _GEN_1399; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1401 = i == 8'hc6 ? _GEN_1400 : _GEN_1399; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1402 = io_inputBit ? 1'h0 : _GEN_1401; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1403 = i == 8'hc6 ? _GEN_1402 : _GEN_1401; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1404 = ~io_inputBit ? 1'h0 : _GEN_1403; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1405 = i == 8'hc7 ? _GEN_1404 : _GEN_1403; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1406 = io_inputBit | _GEN_1405; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1407 = i == 8'hc7 ? _GEN_1406 : _GEN_1405; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1408 = ~io_inputBit | _GEN_1407; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1409 = i == 8'hc9 ? _GEN_1408 : _GEN_1407; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1410 = io_inputBit ? 1'h0 : _GEN_1409; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1411 = i == 8'hc9 ? _GEN_1410 : _GEN_1409; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1412 = ~io_inputBit ? 1'h0 : _GEN_1411; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1413 = i == 8'hca ? _GEN_1412 : _GEN_1411; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1414 = io_inputBit | _GEN_1413; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1415 = i == 8'hca ? _GEN_1414 : _GEN_1413; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1416 = ~io_inputBit | _GEN_1415; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1417 = i == 8'hcb ? _GEN_1416 : _GEN_1415; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1418 = io_inputBit ? 1'h0 : _GEN_1417; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1419 = i == 8'hcb ? _GEN_1418 : _GEN_1417; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1420 = ~io_inputBit ? 1'h0 : _GEN_1419; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1421 = i == 8'hcd ? _GEN_1420 : _GEN_1419; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1422 = io_inputBit | _GEN_1421; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1423 = i == 8'hcd ? _GEN_1422 : _GEN_1421; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1424 = ~io_inputBit | _GEN_1423; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1425 = i == 8'hce ? _GEN_1424 : _GEN_1423; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1428 = ~io_inputBit ? 1'h0 : _GEN_1037; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1429 = i == 8'h1 ? _GEN_1428 : _GEN_1037; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1430 = io_inputBit ? 1'h0 : _GEN_1429; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1431 = i == 8'h2 ? _GEN_1430 : _GEN_1429; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1432 = ~io_inputBit ? 1'h0 : _GEN_1431; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1433 = i == 8'h4 ? _GEN_1432 : _GEN_1431; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1434 = io_inputBit ? 1'h0 : _GEN_1433; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1435 = i == 8'h5 ? _GEN_1434 : _GEN_1433; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1436 = io_inputBit | _GEN_1435; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1437 = i == 8'h16 ? _GEN_1436 : _GEN_1435; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1438 = ~io_inputBit | _GEN_1437; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1439 = i == 8'h17 ? _GEN_1438 : _GEN_1437; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1440 = ~io_inputBit ? 1'h0 : _GEN_1439; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1441 = i == 8'h2b ? _GEN_1440 : _GEN_1439; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1442 = ~io_inputBit | _GEN_1441; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1443 = i == 8'h30 ? _GEN_1442 : _GEN_1441; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1444 = ~io_inputBit | _GEN_1443; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1445 = i == 8'h62 ? _GEN_1444 : _GEN_1443; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1446 = ~io_inputBit ? 1'h0 : _GEN_1445; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1447 = i == 8'h63 ? _GEN_1446 : _GEN_1445; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1448 = ~io_inputBit | _GEN_1447; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1449 = i == 8'h64 ? _GEN_1448 : _GEN_1447; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1450 = ~io_inputBit ? 1'h0 : _GEN_1449; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1451 = i == 8'h65 ? _GEN_1450 : _GEN_1449; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1452 = ~io_inputBit | _GEN_1451; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1453 = i == 8'h66 ? _GEN_1452 : _GEN_1451; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1454 = ~io_inputBit ? 1'h0 : _GEN_1453; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1455 = i == 8'hb1 ? _GEN_1454 : _GEN_1453; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1456 = io_inputBit | _GEN_1455; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1457 = i == 8'hb1 ? _GEN_1456 : _GEN_1455; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1458 = ~io_inputBit ? 1'h0 : _GEN_1457; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1459 = i == 8'hb2 ? _GEN_1458 : _GEN_1457; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1460 = io_inputBit | _GEN_1459; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1461 = i == 8'hb2 ? _GEN_1460 : _GEN_1459; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1462 = ~io_inputBit | _GEN_1461; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1463 = i == 8'hb3 ? _GEN_1462 : _GEN_1461; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1464 = io_inputBit ? 1'h0 : _GEN_1463; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1465 = i == 8'hb3 ? _GEN_1464 : _GEN_1463; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1466 = ~io_inputBit | _GEN_1465; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1467 = i == 8'hb4 ? _GEN_1466 : _GEN_1465; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1468 = io_inputBit ? 1'h0 : _GEN_1467; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1469 = i == 8'hb4 ? _GEN_1468 : _GEN_1467; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1470 = ~io_inputBit ? 1'h0 : _GEN_1469; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1471 = i == 8'hb5 ? _GEN_1470 : _GEN_1469; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1472 = io_inputBit | _GEN_1471; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1473 = i == 8'hb5 ? _GEN_1472 : _GEN_1471; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1474 = ~io_inputBit ? 1'h0 : _GEN_1473; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1475 = i == 8'hb6 ? _GEN_1474 : _GEN_1473; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1476 = io_inputBit | _GEN_1475; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1477 = i == 8'hb6 ? _GEN_1476 : _GEN_1475; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1478 = ~io_inputBit | _GEN_1477; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1479 = i == 8'hb7 ? _GEN_1478 : _GEN_1477; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1480 = io_inputBit ? 1'h0 : _GEN_1479; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1481 = i == 8'hb7 ? _GEN_1480 : _GEN_1479; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1482 = ~io_inputBit | _GEN_1481; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1483 = i == 8'hb8 ? _GEN_1482 : _GEN_1481; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1484 = io_inputBit ? 1'h0 : _GEN_1483; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1485 = i == 8'hb8 ? _GEN_1484 : _GEN_1483; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1486 = ~io_inputBit ? 1'h0 : _GEN_1485; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1487 = i == 8'hb9 ? _GEN_1486 : _GEN_1485; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1488 = io_inputBit | _GEN_1487; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1489 = i == 8'hb9 ? _GEN_1488 : _GEN_1487; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1490 = ~io_inputBit ? 1'h0 : _GEN_1489; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1491 = i == 8'hba ? _GEN_1490 : _GEN_1489; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1492 = io_inputBit | _GEN_1491; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1493 = i == 8'hba ? _GEN_1492 : _GEN_1491; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1494 = ~io_inputBit ? 1'h0 : _GEN_1493; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1495 = i == 8'hc6 ? _GEN_1494 : _GEN_1493; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1496 = io_inputBit | _GEN_1495; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1497 = i == 8'hc6 ? _GEN_1496 : _GEN_1495; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1498 = ~io_inputBit | _GEN_1497; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1499 = i == 8'hc8 ? _GEN_1498 : _GEN_1497; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1500 = io_inputBit ? 1'h0 : _GEN_1499; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1501 = i == 8'hc8 ? _GEN_1500 : _GEN_1499; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1502 = ~io_inputBit ? 1'h0 : _GEN_1501; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1503 = i == 8'hca ? _GEN_1502 : _GEN_1501; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1504 = io_inputBit | _GEN_1503; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1505 = i == 8'hca ? _GEN_1504 : _GEN_1503; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1506 = ~io_inputBit | _GEN_1505; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1507 = i == 8'hcc ? _GEN_1506 : _GEN_1505; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1508 = io_inputBit ? 1'h0 : _GEN_1507; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1509 = i == 8'hcc ? _GEN_1508 : _GEN_1507; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1510 = ~io_inputBit ? 1'h0 : _GEN_1509; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1511 = i == 8'hce ? _GEN_1510 : _GEN_1509; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1512 = io_inputBit | _GEN_1511; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1514 = ~io_inputBit ? 1'h0 : _GEN_1113; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1515 = i == 8'h1 ? _GEN_1514 : _GEN_1113; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1516 = io_inputBit ? 1'h0 : _GEN_1515; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1517 = i == 8'h2 ? _GEN_1516 : _GEN_1515; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1518 = ~io_inputBit ? 1'h0 : _GEN_1517; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1519 = i == 8'h4 ? _GEN_1518 : _GEN_1517; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1520 = io_inputBit ? 1'h0 : _GEN_1519; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1521 = i == 8'h5 ? _GEN_1520 : _GEN_1519; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1522 = io_inputBit ? 1'h0 : _GEN_1521; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1523 = i == 8'h16 ? _GEN_1522 : _GEN_1521; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1524 = ~io_inputBit ? 1'h0 : _GEN_1523; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1525 = i == 8'h17 ? _GEN_1524 : _GEN_1523; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1526 = ~io_inputBit ? 1'h0 : _GEN_1525; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1527 = i == 8'h2b ? _GEN_1526 : _GEN_1525; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1528 = ~io_inputBit ? 1'h0 : _GEN_1527; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1529 = i == 8'h30 ? _GEN_1528 : _GEN_1527; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1530 = ~io_inputBit ? 1'h0 : _GEN_1529; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1531 = i == 8'h58 ? _GEN_1530 : _GEN_1529; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1532 = io_inputBit | _GEN_1531; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1533 = i == 8'h58 ? _GEN_1532 : _GEN_1531; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1534 = ~io_inputBit ? 1'h0 : _GEN_1533; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1535 = i == 8'h59 ? _GEN_1534 : _GEN_1533; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1536 = io_inputBit | _GEN_1535; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1537 = i == 8'h59 ? _GEN_1536 : _GEN_1535; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1538 = ~io_inputBit ? 1'h0 : _GEN_1537; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1539 = i == 8'h5a ? _GEN_1538 : _GEN_1537; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1540 = io_inputBit | _GEN_1539; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1541 = i == 8'h5a ? _GEN_1540 : _GEN_1539; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1542 = ~io_inputBit ? 1'h0 : _GEN_1541; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1543 = i == 8'h5b ? _GEN_1542 : _GEN_1541; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1544 = io_inputBit | _GEN_1543; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1545 = i == 8'h5b ? _GEN_1544 : _GEN_1543; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1546 = ~io_inputBit ? 1'h0 : _GEN_1545; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1547 = i == 8'h5c ? _GEN_1546 : _GEN_1545; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1548 = io_inputBit | _GEN_1547; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1549 = i == 8'h5c ? _GEN_1548 : _GEN_1547; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1550 = ~io_inputBit ? 1'h0 : _GEN_1549; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1551 = i == 8'hc5 ? _GEN_1550 : _GEN_1549; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1552 = io_inputBit | _GEN_1551; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1553 = i == 8'hc5 ? _GEN_1552 : _GEN_1551; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1554 = ~io_inputBit | _GEN_1553; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1555 = i == 8'hc6 ? _GEN_1554 : _GEN_1553; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1556 = io_inputBit ? 1'h0 : _GEN_1555; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1557 = i == 8'hc6 ? _GEN_1556 : _GEN_1555; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1558 = ~io_inputBit ? 1'h0 : _GEN_1557; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1559 = i == 8'hc7 ? _GEN_1558 : _GEN_1557; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1560 = io_inputBit | _GEN_1559; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1561 = i == 8'hc7 ? _GEN_1560 : _GEN_1559; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1562 = ~io_inputBit | _GEN_1561; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1563 = i == 8'hc8 ? _GEN_1562 : _GEN_1561; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1564 = io_inputBit ? 1'h0 : _GEN_1563; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1565 = i == 8'hc8 ? _GEN_1564 : _GEN_1563; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1566 = ~io_inputBit ? 1'h0 : _GEN_1565; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1567 = i == 8'hc9 ? _GEN_1566 : _GEN_1565; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1568 = io_inputBit | _GEN_1567; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1569 = i == 8'hc9 ? _GEN_1568 : _GEN_1567; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1570 = ~io_inputBit | _GEN_1569; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1571 = i == 8'hca ? _GEN_1570 : _GEN_1569; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1572 = io_inputBit ? 1'h0 : _GEN_1571; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1573 = i == 8'hca ? _GEN_1572 : _GEN_1571; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1574 = ~io_inputBit ? 1'h0 : _GEN_1573; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1575 = i == 8'hcb ? _GEN_1574 : _GEN_1573; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1576 = io_inputBit | _GEN_1575; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1577 = i == 8'hcb ? _GEN_1576 : _GEN_1575; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1578 = ~io_inputBit | _GEN_1577; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1579 = i == 8'hcc ? _GEN_1578 : _GEN_1577; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1580 = io_inputBit ? 1'h0 : _GEN_1579; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1581 = i == 8'hcc ? _GEN_1580 : _GEN_1579; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1582 = ~io_inputBit ? 1'h0 : _GEN_1581; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1583 = i == 8'hcd ? _GEN_1582 : _GEN_1581; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1584 = io_inputBit | _GEN_1583; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1585 = i == 8'hcd ? _GEN_1584 : _GEN_1583; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1586 = ~io_inputBit | _GEN_1585; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1587 = i == 8'hce ? _GEN_1586 : _GEN_1585; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1590 = ~io_inputBit ? 1'h0 : _GEN_1209; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1591 = i == 8'h1 ? _GEN_1590 : _GEN_1209; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1592 = io_inputBit ? 1'h0 : _GEN_1591; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1593 = i == 8'h2 ? _GEN_1592 : _GEN_1591; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1594 = ~io_inputBit ? 1'h0 : _GEN_1593; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1595 = i == 8'h4 ? _GEN_1594 : _GEN_1593; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1596 = io_inputBit ? 1'h0 : _GEN_1595; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1597 = i == 8'h5 ? _GEN_1596 : _GEN_1595; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1598 = io_inputBit ? 1'h0 : _GEN_1597; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1599 = i == 8'h16 ? _GEN_1598 : _GEN_1597; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1600 = ~io_inputBit ? 1'h0 : _GEN_1599; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1601 = i == 8'h17 ? _GEN_1600 : _GEN_1599; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1602 = ~io_inputBit ? 1'h0 : _GEN_1601; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1603 = i == 8'h2b ? _GEN_1602 : _GEN_1601; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1604 = ~io_inputBit ? 1'h0 : _GEN_1603; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1605 = i == 8'h30 ? _GEN_1604 : _GEN_1603; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1606 = ~io_inputBit ? 1'h0 : _GEN_1605; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1607 = i == 8'hb1 ? _GEN_1606 : _GEN_1605; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1608 = io_inputBit | _GEN_1607; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1609 = i == 8'hb1 ? _GEN_1608 : _GEN_1607; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1610 = ~io_inputBit ? 1'h0 : _GEN_1609; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1611 = i == 8'hb2 ? _GEN_1610 : _GEN_1609; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1612 = io_inputBit | _GEN_1611; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1613 = i == 8'hb2 ? _GEN_1612 : _GEN_1611; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1614 = ~io_inputBit ? 1'h0 : _GEN_1613; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1615 = i == 8'hb3 ? _GEN_1614 : _GEN_1613; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1616 = io_inputBit | _GEN_1615; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1617 = i == 8'hb3 ? _GEN_1616 : _GEN_1615; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1618 = ~io_inputBit ? 1'h0 : _GEN_1617; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1619 = i == 8'hb4 ? _GEN_1618 : _GEN_1617; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1620 = io_inputBit | _GEN_1619; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1621 = i == 8'hb4 ? _GEN_1620 : _GEN_1619; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1622 = ~io_inputBit ? 1'h0 : _GEN_1621; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1623 = i == 8'hb5 ? _GEN_1622 : _GEN_1621; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1624 = io_inputBit | _GEN_1623; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1625 = i == 8'hb5 ? _GEN_1624 : _GEN_1623; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1626 = ~io_inputBit ? 1'h0 : _GEN_1625; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1627 = i == 8'hb6 ? _GEN_1626 : _GEN_1625; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1628 = io_inputBit | _GEN_1627; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1629 = i == 8'hb6 ? _GEN_1628 : _GEN_1627; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1630 = ~io_inputBit ? 1'h0 : _GEN_1629; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1631 = i == 8'hb7 ? _GEN_1630 : _GEN_1629; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1632 = io_inputBit | _GEN_1631; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1633 = i == 8'hb7 ? _GEN_1632 : _GEN_1631; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1634 = ~io_inputBit ? 1'h0 : _GEN_1633; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1635 = i == 8'hb8 ? _GEN_1634 : _GEN_1633; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1636 = io_inputBit | _GEN_1635; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1637 = i == 8'hb8 ? _GEN_1636 : _GEN_1635; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1638 = ~io_inputBit ? 1'h0 : _GEN_1637; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1639 = i == 8'hb9 ? _GEN_1638 : _GEN_1637; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1640 = io_inputBit | _GEN_1639; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1641 = i == 8'hb9 ? _GEN_1640 : _GEN_1639; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1642 = ~io_inputBit ? 1'h0 : _GEN_1641; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1643 = i == 8'hba ? _GEN_1642 : _GEN_1641; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1644 = io_inputBit | _GEN_1643; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1645 = i == 8'hba ? _GEN_1644 : _GEN_1643; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1646 = ~io_inputBit ? 1'h0 : _GEN_1645; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1647 = i == 8'hc5 ? _GEN_1646 : _GEN_1645; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1648 = io_inputBit | _GEN_1647; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1649 = i == 8'hc5 ? _GEN_1648 : _GEN_1647; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1650 = ~io_inputBit ? 1'h0 : _GEN_1649; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1651 = i == 8'hc6 ? _GEN_1650 : _GEN_1649; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1652 = io_inputBit | _GEN_1651; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1653 = i == 8'hc6 ? _GEN_1652 : _GEN_1651; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1654 = ~io_inputBit ? 1'h0 : _GEN_1653; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1655 = i == 8'hc7 ? _GEN_1654 : _GEN_1653; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1656 = io_inputBit | _GEN_1655; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1657 = i == 8'hc7 ? _GEN_1656 : _GEN_1655; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1658 = ~io_inputBit ? 1'h0 : _GEN_1657; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1659 = i == 8'hc8 ? _GEN_1658 : _GEN_1657; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1660 = io_inputBit | _GEN_1659; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1661 = i == 8'hc8 ? _GEN_1660 : _GEN_1659; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1662 = ~io_inputBit ? 1'h0 : _GEN_1661; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1663 = i == 8'hc9 ? _GEN_1662 : _GEN_1661; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1664 = io_inputBit | _GEN_1663; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1665 = i == 8'hc9 ? _GEN_1664 : _GEN_1663; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1666 = ~io_inputBit ? 1'h0 : _GEN_1665; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1667 = i == 8'hca ? _GEN_1666 : _GEN_1665; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1668 = io_inputBit | _GEN_1667; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1669 = i == 8'hca ? _GEN_1668 : _GEN_1667; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1670 = ~io_inputBit ? 1'h0 : _GEN_1669; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1671 = i == 8'hcb ? _GEN_1670 : _GEN_1669; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1672 = io_inputBit | _GEN_1671; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1673 = i == 8'hcb ? _GEN_1672 : _GEN_1671; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1674 = ~io_inputBit ? 1'h0 : _GEN_1673; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1675 = i == 8'hcc ? _GEN_1674 : _GEN_1673; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1676 = io_inputBit | _GEN_1675; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1677 = i == 8'hcc ? _GEN_1676 : _GEN_1675; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1678 = ~io_inputBit ? 1'h0 : _GEN_1677; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1679 = i == 8'hcd ? _GEN_1678 : _GEN_1677; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1680 = io_inputBit | _GEN_1679; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1681 = i == 8'hcd ? _GEN_1680 : _GEN_1679; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1682 = ~io_inputBit ? 1'h0 : _GEN_1681; // @[lut_mem_online.scala 236:46 238:32]
  wire  _GEN_1683 = i == 8'hce ? _GEN_1682 : _GEN_1681; // @[lut_mem_online.scala 234:34]
  wire  _GEN_1684 = io_inputBit | _GEN_1683; // @[lut_mem_online.scala 236:46 238:32]
  wire  _T_1689 = counter < 4'hf; // @[lut_mem_online.scala 248:22]
  wire  _T_1691 = counter >= 4'h8; // @[lut_mem_online.scala 256:30]
  wire [3:0] _outResult_T_1 = counter - 4'h8; // @[lut_mem_online.scala 258:41]
  wire  _GEN_1694 = 3'h1 == _outResult_T_1[2:0] ? buffer_1 : buffer_0; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_1695 = 3'h2 == _outResult_T_1[2:0] ? buffer_2 : _GEN_1694; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_1696 = 3'h3 == _outResult_T_1[2:0] ? buffer_3 : _GEN_1695; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_1697 = 3'h4 == _outResult_T_1[2:0] ? buffer_4 : _GEN_1696; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_1698 = 3'h5 == _outResult_T_1[2:0] ? buffer_5 : _GEN_1697; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_1699 = 3'h6 == _outResult_T_1[2:0] ? buffer_6 : _GEN_1698; // @[lut_mem_online.scala 258:{23,23}]
  wire  _GEN_1700 = 3'h7 == _outResult_T_1[2:0] ? 1'h0 : _GEN_1699; // @[lut_mem_online.scala 258:{23,23}]
  wire  _T_1695 = ~reset; // @[lut_mem_online.scala 260:21]
  wire  _GEN_1702 = counter >= 4'h8 ? _GEN_1700 : outResult; // @[lut_mem_online.scala 256:42 258:23 214:26]
  wire  _GEN_1704 = _T_2 ? 1'h0 : _GEN_1702; // @[lut_mem_online.scala 253:35 255:23]
  wire  _T_1696 = i < 8'h7f; // @[lut_mem_online.scala 271:18]
  wire [9:0] _i_T = 2'h2 * i; // @[lut_mem_online.scala 281:24]
  wire [9:0] _i_T_2 = _i_T + 10'h1; // @[lut_mem_online.scala 281:28]
  wire [9:0] _i_T_5 = _i_T + 10'h2; // @[lut_mem_online.scala 283:28]
  wire [9:0] _GEN_1705 = io_inputBit ? _i_T_5 : {{2'd0}, i}; // @[lut_mem_online.scala 282:45 283:17 205:18]
  wire [9:0] _GEN_1706 = _T_10 ? _i_T_2 : _GEN_1705; // @[lut_mem_online.scala 280:39 281:17]
  wire  _T_1701 = i < 8'hff; // @[lut_mem_online.scala 286:24]
  wire [7:0] _GEN_1707 = i < 8'hff ? 8'hff : i; // @[lut_mem_online.scala 286:63 294:15 205:18]
  wire [9:0] _GEN_1708 = i < 8'h7f ? _GEN_1706 : {{2'd0}, _GEN_1707}; // @[lut_mem_online.scala 271:61]
  wire [3:0] _counter_T_1 = counter + 4'h1; // @[lut_mem_online.scala 297:30]
  wire  _GEN_1710 = counter < 4'hf & _GEN_1704; // @[lut_mem_online.scala 248:52 300:21]
  wire [9:0] _GEN_1711 = counter < 4'hf ? _GEN_1708 : {{2'd0}, i}; // @[lut_mem_online.scala 205:18 248:52]
  wire  _GEN_1734 = io_start & _GEN_1710; // @[lut_mem_online.scala 219:29 323:15]
  wire [9:0] _GEN_1735 = io_start ? _GEN_1711 : 10'h0; // @[lut_mem_online.scala 219:29 321:7]
  wire [9:0] _GEN_1738 = reset ? 10'h0 : _GEN_1735; // @[lut_mem_online.scala 205:{18,18}]
  wire  _GEN_1739 = io_start & _T_1689; // @[lut_mem_online.scala 260:21]
  assign io_outResult = outResult; // @[lut_mem_online.scala 330:16]
  always @(posedge clock) begin
    i <= _GEN_1738[7:0]; // @[lut_mem_online.scala 205:{18,18}]
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hb7) begin // @[lut_mem_online.scala 234:34]
          buffer_0 <= _GEN_1236;
        end else if (i == 8'hb7) begin // @[lut_mem_online.scala 234:34]
          buffer_0 <= _GEN_1234;
        end else begin
          buffer_0 <= _GEN_1233;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hc5) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_1 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_1 <= _GEN_1283;
          end
        end else begin
          buffer_1 <= _GEN_1283;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hcd) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_2 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_2 <= _GEN_1345;
          end
        end else begin
          buffer_2 <= _GEN_1345;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hce) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_3 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_3 <= _GEN_1425;
          end
        end else begin
          buffer_3 <= _GEN_1425;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hce) begin // @[lut_mem_online.scala 234:34]
          buffer_4 <= _GEN_1512;
        end else if (i == 8'hce) begin // @[lut_mem_online.scala 234:34]
          buffer_4 <= _GEN_1510;
        end else begin
          buffer_4 <= _GEN_1509;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hce) begin // @[lut_mem_online.scala 234:34]
          if (io_inputBit) begin // @[lut_mem_online.scala 236:46]
            buffer_5 <= 1'h0; // @[lut_mem_online.scala 238:32]
          end else begin
            buffer_5 <= _GEN_1587;
          end
        end else begin
          buffer_5 <= _GEN_1587;
        end
      end
    end
    if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'h8) begin // @[lut_mem_online.scala 231:36]
        if (i == 8'hce) begin // @[lut_mem_online.scala 234:34]
          buffer_6 <= _GEN_1684;
        end else if (i == 8'hce) begin // @[lut_mem_online.scala 234:34]
          buffer_6 <= _GEN_1682;
        end else begin
          buffer_6 <= _GEN_1681;
        end
      end
    end
    if (reset) begin // @[lut_mem_online.scala 211:24]
      counter <= 4'h0; // @[lut_mem_online.scala 211:24]
    end else if (io_start) begin // @[lut_mem_online.scala 219:29]
      if (counter < 4'hf) begin // @[lut_mem_online.scala 248:52]
        counter <= _counter_T_1; // @[lut_mem_online.scala 297:19]
      end
    end else begin
      counter <= 4'h0; // @[lut_mem_online.scala 322:13]
    end
    if (reset) begin // @[lut_mem_online.scala 214:26]
      outResult <= 1'h0; // @[lut_mem_online.scala 214:26]
    end else begin
      outResult <= _GEN_1734;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & _T_1689 & ~_T_2 & _T_1691 & ~reset) begin
          $fwrite(32'h80000002,"debug, set buffer to output buffer(%d), counter = %d\n",_outResult_T_1,counter); // @[lut_mem_online.scala 260:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1739 & _T_1696 & _T_1695) begin
          $fwrite(32'h80000002,"debug, state transition 1: %d\n",i); // @[lut_mem_online.scala 274:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1739 & ~_T_1696 & _T_1701 & _T_1695) begin
          $fwrite(32'h80000002,"debug, state transition 2: %d\n",i); // @[lut_mem_online.scala 289:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
