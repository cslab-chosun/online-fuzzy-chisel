module RegularFuzzification(
  input        clock,
  input        reset,
  input        io_start,
  input  [9:0] io_inputs_0,
  input  [9:0] io_inputs_1,
  output       io_outResultValid,
  output [2:0] io_outResult
);
  wire  regMaxVec_0_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_0_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_0_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_1_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_1_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_inputs_5; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_1_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_2_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_2_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_2_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_3_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_3_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_inputs_5; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_3_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_4_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_4_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] regMaxVec_4_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  outResult_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  outResult_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [2:0] outResult_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  reg [2:0] regLutResultsVec_0; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_1; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_2; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_3; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regLutResultsVec_4; // @[regular_fuzzification.scala 125:29]
  reg [2:0] regMinVec_0; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_1; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_2; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_3; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_4; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_5; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_6; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_7; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_8; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_9; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_10; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_11; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_12; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_13; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_14; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_15; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_16; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_17; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_18; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_19; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_20; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_21; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_22; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_23; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMinVec_24; // @[regular_fuzzification.scala 144:22]
  reg [2:0] regMaxVec_0; // @[regular_fuzzification.scala 158:22]
  reg [2:0] regMaxVec_1; // @[regular_fuzzification.scala 158:22]
  reg [2:0] regMaxVec_2; // @[regular_fuzzification.scala 158:22]
  reg [2:0] regMaxVec_3; // @[regular_fuzzification.scala 158:22]
  reg [2:0] regMaxVec_4; // @[regular_fuzzification.scala 158:22]
  wire [6:0] _GEN_21 = 8'h15 == io_inputs_0[7:0] ? 7'h5f : 7'h64; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_22 = 8'h16 == io_inputs_0[7:0] ? 7'h5a : _GEN_21; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_23 = 8'h17 == io_inputs_0[7:0] ? 7'h55 : _GEN_22; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_24 = 8'h18 == io_inputs_0[7:0] ? 7'h50 : _GEN_23; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_25 = 8'h19 == io_inputs_0[7:0] ? 7'h4b : _GEN_24; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_26 = 8'h1a == io_inputs_0[7:0] ? 7'h46 : _GEN_25; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_27 = 8'h1b == io_inputs_0[7:0] ? 7'h41 : _GEN_26; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_28 = 8'h1c == io_inputs_0[7:0] ? 7'h3c : _GEN_27; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_29 = 8'h1d == io_inputs_0[7:0] ? 7'h37 : _GEN_28; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_30 = 8'h1e == io_inputs_0[7:0] ? 7'h32 : _GEN_29; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_31 = 8'h1f == io_inputs_0[7:0] ? 7'h2d : _GEN_30; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_32 = 8'h20 == io_inputs_0[7:0] ? 7'h28 : _GEN_31; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_33 = 8'h21 == io_inputs_0[7:0] ? 7'h23 : _GEN_32; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_34 = 8'h22 == io_inputs_0[7:0] ? 7'h1e : _GEN_33; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_35 = 8'h23 == io_inputs_0[7:0] ? 7'h19 : _GEN_34; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_36 = 8'h24 == io_inputs_0[7:0] ? 7'h14 : _GEN_35; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_37 = 8'h25 == io_inputs_0[7:0] ? 7'hf : _GEN_36; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_38 = 8'h26 == io_inputs_0[7:0] ? 7'ha : _GEN_37; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_39 = 8'h27 == io_inputs_0[7:0] ? 7'h5 : _GEN_38; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_40 = 8'h28 == io_inputs_0[7:0] ? 7'h0 : _GEN_39; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_41 = 8'h29 == io_inputs_0[7:0] ? 7'h0 : _GEN_40; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_42 = 8'h2a == io_inputs_0[7:0] ? 7'h0 : _GEN_41; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_43 = 8'h2b == io_inputs_0[7:0] ? 7'h0 : _GEN_42; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_44 = 8'h2c == io_inputs_0[7:0] ? 7'h0 : _GEN_43; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_45 = 8'h2d == io_inputs_0[7:0] ? 7'h0 : _GEN_44; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_46 = 8'h2e == io_inputs_0[7:0] ? 7'h0 : _GEN_45; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_47 = 8'h2f == io_inputs_0[7:0] ? 7'h0 : _GEN_46; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_48 = 8'h30 == io_inputs_0[7:0] ? 7'h0 : _GEN_47; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_49 = 8'h31 == io_inputs_0[7:0] ? 7'h0 : _GEN_48; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_50 = 8'h32 == io_inputs_0[7:0] ? 7'h0 : _GEN_49; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_51 = 8'h33 == io_inputs_0[7:0] ? 7'h0 : _GEN_50; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_52 = 8'h34 == io_inputs_0[7:0] ? 7'h0 : _GEN_51; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_53 = 8'h35 == io_inputs_0[7:0] ? 7'h0 : _GEN_52; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_54 = 8'h36 == io_inputs_0[7:0] ? 7'h0 : _GEN_53; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_55 = 8'h37 == io_inputs_0[7:0] ? 7'h0 : _GEN_54; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_56 = 8'h38 == io_inputs_0[7:0] ? 7'h0 : _GEN_55; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_57 = 8'h39 == io_inputs_0[7:0] ? 7'h0 : _GEN_56; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_58 = 8'h3a == io_inputs_0[7:0] ? 7'h0 : _GEN_57; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_59 = 8'h3b == io_inputs_0[7:0] ? 7'h0 : _GEN_58; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_60 = 8'h3c == io_inputs_0[7:0] ? 7'h0 : _GEN_59; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_61 = 8'h3d == io_inputs_0[7:0] ? 7'h0 : _GEN_60; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_62 = 8'h3e == io_inputs_0[7:0] ? 7'h0 : _GEN_61; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_63 = 8'h3f == io_inputs_0[7:0] ? 7'h0 : _GEN_62; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_64 = 8'h40 == io_inputs_0[7:0] ? 7'h0 : _GEN_63; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_65 = 8'h41 == io_inputs_0[7:0] ? 7'h0 : _GEN_64; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_66 = 8'h42 == io_inputs_0[7:0] ? 7'h0 : _GEN_65; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_67 = 8'h43 == io_inputs_0[7:0] ? 7'h0 : _GEN_66; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_68 = 8'h44 == io_inputs_0[7:0] ? 7'h0 : _GEN_67; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_69 = 8'h45 == io_inputs_0[7:0] ? 7'h0 : _GEN_68; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_70 = 8'h46 == io_inputs_0[7:0] ? 7'h0 : _GEN_69; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_71 = 8'h47 == io_inputs_0[7:0] ? 7'h0 : _GEN_70; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_72 = 8'h48 == io_inputs_0[7:0] ? 7'h0 : _GEN_71; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_73 = 8'h49 == io_inputs_0[7:0] ? 7'h0 : _GEN_72; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_74 = 8'h4a == io_inputs_0[7:0] ? 7'h0 : _GEN_73; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_75 = 8'h4b == io_inputs_0[7:0] ? 7'h0 : _GEN_74; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_76 = 8'h4c == io_inputs_0[7:0] ? 7'h0 : _GEN_75; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_77 = 8'h4d == io_inputs_0[7:0] ? 7'h0 : _GEN_76; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_78 = 8'h4e == io_inputs_0[7:0] ? 7'h0 : _GEN_77; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_79 = 8'h4f == io_inputs_0[7:0] ? 7'h0 : _GEN_78; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_80 = 8'h50 == io_inputs_0[7:0] ? 7'h0 : _GEN_79; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_81 = 8'h51 == io_inputs_0[7:0] ? 7'h0 : _GEN_80; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_82 = 8'h52 == io_inputs_0[7:0] ? 7'h0 : _GEN_81; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_83 = 8'h53 == io_inputs_0[7:0] ? 7'h0 : _GEN_82; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_84 = 8'h54 == io_inputs_0[7:0] ? 7'h0 : _GEN_83; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_85 = 8'h55 == io_inputs_0[7:0] ? 7'h0 : _GEN_84; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_86 = 8'h56 == io_inputs_0[7:0] ? 7'h0 : _GEN_85; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_87 = 8'h57 == io_inputs_0[7:0] ? 7'h0 : _GEN_86; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_88 = 8'h58 == io_inputs_0[7:0] ? 7'h0 : _GEN_87; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_89 = 8'h59 == io_inputs_0[7:0] ? 7'h0 : _GEN_88; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_90 = 8'h5a == io_inputs_0[7:0] ? 7'h0 : _GEN_89; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_91 = 8'h5b == io_inputs_0[7:0] ? 7'h0 : _GEN_90; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_92 = 8'h5c == io_inputs_0[7:0] ? 7'h0 : _GEN_91; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_93 = 8'h5d == io_inputs_0[7:0] ? 7'h0 : _GEN_92; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_94 = 8'h5e == io_inputs_0[7:0] ? 7'h0 : _GEN_93; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_95 = 8'h5f == io_inputs_0[7:0] ? 7'h0 : _GEN_94; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_96 = 8'h60 == io_inputs_0[7:0] ? 7'h0 : _GEN_95; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_97 = 8'h61 == io_inputs_0[7:0] ? 7'h0 : _GEN_96; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_98 = 8'h62 == io_inputs_0[7:0] ? 7'h0 : _GEN_97; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_99 = 8'h63 == io_inputs_0[7:0] ? 7'h0 : _GEN_98; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_100 = 8'h64 == io_inputs_0[7:0] ? 7'h0 : _GEN_99; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_101 = 8'h65 == io_inputs_0[7:0] ? 7'h0 : _GEN_100; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_102 = 8'h66 == io_inputs_0[7:0] ? 7'h0 : _GEN_101; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_103 = 8'h67 == io_inputs_0[7:0] ? 7'h0 : _GEN_102; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_104 = 8'h68 == io_inputs_0[7:0] ? 7'h0 : _GEN_103; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_105 = 8'h69 == io_inputs_0[7:0] ? 7'h0 : _GEN_104; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_106 = 8'h6a == io_inputs_0[7:0] ? 7'h0 : _GEN_105; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_107 = 8'h6b == io_inputs_0[7:0] ? 7'h0 : _GEN_106; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_108 = 8'h6c == io_inputs_0[7:0] ? 7'h0 : _GEN_107; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_109 = 8'h6d == io_inputs_0[7:0] ? 7'h0 : _GEN_108; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_110 = 8'h6e == io_inputs_0[7:0] ? 7'h0 : _GEN_109; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_111 = 8'h6f == io_inputs_0[7:0] ? 7'h0 : _GEN_110; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_112 = 8'h70 == io_inputs_0[7:0] ? 7'h0 : _GEN_111; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_113 = 8'h71 == io_inputs_0[7:0] ? 7'h0 : _GEN_112; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_114 = 8'h72 == io_inputs_0[7:0] ? 7'h0 : _GEN_113; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_115 = 8'h73 == io_inputs_0[7:0] ? 7'h0 : _GEN_114; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_116 = 8'h74 == io_inputs_0[7:0] ? 7'h0 : _GEN_115; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_117 = 8'h75 == io_inputs_0[7:0] ? 7'h0 : _GEN_116; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_118 = 8'h76 == io_inputs_0[7:0] ? 7'h0 : _GEN_117; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_119 = 8'h77 == io_inputs_0[7:0] ? 7'h0 : _GEN_118; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_120 = 8'h78 == io_inputs_0[7:0] ? 7'h0 : _GEN_119; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_121 = 8'h79 == io_inputs_0[7:0] ? 7'h0 : _GEN_120; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_122 = 8'h7a == io_inputs_0[7:0] ? 7'h0 : _GEN_121; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_123 = 8'h7b == io_inputs_0[7:0] ? 7'h0 : _GEN_122; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_124 = 8'h7c == io_inputs_0[7:0] ? 7'h0 : _GEN_123; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_125 = 8'h7d == io_inputs_0[7:0] ? 7'h0 : _GEN_124; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_126 = 8'h7e == io_inputs_0[7:0] ? 7'h0 : _GEN_125; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_127 = 8'h7f == io_inputs_0[7:0] ? 7'h0 : _GEN_126; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_128 = 8'h80 == io_inputs_0[7:0] ? 7'h0 : _GEN_127; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_129 = 8'h81 == io_inputs_0[7:0] ? 7'h0 : _GEN_128; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_130 = 8'h82 == io_inputs_0[7:0] ? 7'h0 : _GEN_129; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_131 = 8'h83 == io_inputs_0[7:0] ? 7'h0 : _GEN_130; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_132 = 8'h84 == io_inputs_0[7:0] ? 7'h0 : _GEN_131; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_133 = 8'h85 == io_inputs_0[7:0] ? 7'h0 : _GEN_132; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_134 = 8'h86 == io_inputs_0[7:0] ? 7'h0 : _GEN_133; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_135 = 8'h87 == io_inputs_0[7:0] ? 7'h0 : _GEN_134; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_136 = 8'h88 == io_inputs_0[7:0] ? 7'h0 : _GEN_135; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_137 = 8'h89 == io_inputs_0[7:0] ? 7'h0 : _GEN_136; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_138 = 8'h8a == io_inputs_0[7:0] ? 7'h0 : _GEN_137; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_139 = 8'h8b == io_inputs_0[7:0] ? 7'h0 : _GEN_138; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_140 = 8'h8c == io_inputs_0[7:0] ? 7'h0 : _GEN_139; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_141 = 8'h8d == io_inputs_0[7:0] ? 7'h0 : _GEN_140; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_142 = 8'h8e == io_inputs_0[7:0] ? 7'h0 : _GEN_141; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_143 = 8'h8f == io_inputs_0[7:0] ? 7'h0 : _GEN_142; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_144 = 8'h90 == io_inputs_0[7:0] ? 7'h0 : _GEN_143; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_145 = 8'h91 == io_inputs_0[7:0] ? 7'h0 : _GEN_144; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_146 = 8'h92 == io_inputs_0[7:0] ? 7'h0 : _GEN_145; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_147 = 8'h93 == io_inputs_0[7:0] ? 7'h0 : _GEN_146; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_148 = 8'h94 == io_inputs_0[7:0] ? 7'h0 : _GEN_147; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_149 = 8'h95 == io_inputs_0[7:0] ? 7'h0 : _GEN_148; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_150 = 8'h96 == io_inputs_0[7:0] ? 7'h0 : _GEN_149; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_151 = 8'h97 == io_inputs_0[7:0] ? 7'h0 : _GEN_150; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_152 = 8'h98 == io_inputs_0[7:0] ? 7'h0 : _GEN_151; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_153 = 8'h99 == io_inputs_0[7:0] ? 7'h0 : _GEN_152; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_154 = 8'h9a == io_inputs_0[7:0] ? 7'h0 : _GEN_153; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_155 = 8'h9b == io_inputs_0[7:0] ? 7'h0 : _GEN_154; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_156 = 8'h9c == io_inputs_0[7:0] ? 7'h0 : _GEN_155; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_157 = 8'h9d == io_inputs_0[7:0] ? 7'h0 : _GEN_156; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_158 = 8'h9e == io_inputs_0[7:0] ? 7'h0 : _GEN_157; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_159 = 8'h9f == io_inputs_0[7:0] ? 7'h0 : _GEN_158; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_160 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_159; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_161 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_160; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_162 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_161; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_163 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_162; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_164 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_163; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_165 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_164; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_166 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_165; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_167 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_166; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_168 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_167; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_169 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_168; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_170 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_169; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_171 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_170; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_172 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_171; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_173 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_172; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_174 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_173; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_175 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_174; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_176 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_175; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_177 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_176; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_178 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_177; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_179 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_178; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_180 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_179; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_181 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_180; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_182 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_181; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_183 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_182; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_184 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_183; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_185 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_184; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_186 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_185; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_187 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_186; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_188 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_187; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_189 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_188; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_190 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_189; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_191 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_190; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_192 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_191; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_193 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_192; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_194 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_193; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_195 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_194; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_196 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_195; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_197 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_196; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_198 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_197; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_199 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_198; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_200 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_199; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_201 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_200; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_202 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_201; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_203 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_202; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_204 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_203; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_205 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_204; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_206 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_205; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_207 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_206; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_208 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_207; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_209 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_208; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_210 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_209; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_211 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_210; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_212 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_211; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_213 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_212; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_214 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_213; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_215 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_214; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_216 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_215; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_217 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_216; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_218 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_217; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_219 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_218; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_220 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_219; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_221 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_220; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_222 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_221; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_223 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_222; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_224 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_223; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_225 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_224; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_226 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_225; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_227 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_226; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_228 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_227; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_229 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_228; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_230 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_229; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_231 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_230; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_232 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_231; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_233 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_232; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_234 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_233; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_235 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_234; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_236 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_235; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_237 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_236; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_238 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_237; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_239 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_238; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_240 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_239; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_241 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_240; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_242 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_241; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_243 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_242; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_244 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_243; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_245 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_244; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_246 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_245; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_247 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_246; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_248 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_247; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_249 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_248; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_250 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_249; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_251 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_250; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_252 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_251; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_253 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_252; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_254 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_253; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_255 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_254; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_277 = 8'h15 == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_278 = 8'h16 == io_inputs_0[7:0] ? 7'ha : _GEN_277; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_279 = 8'h17 == io_inputs_0[7:0] ? 7'hf : _GEN_278; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_280 = 8'h18 == io_inputs_0[7:0] ? 7'h14 : _GEN_279; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_281 = 8'h19 == io_inputs_0[7:0] ? 7'h19 : _GEN_280; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_282 = 8'h1a == io_inputs_0[7:0] ? 7'h1e : _GEN_281; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_283 = 8'h1b == io_inputs_0[7:0] ? 7'h23 : _GEN_282; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_284 = 8'h1c == io_inputs_0[7:0] ? 7'h28 : _GEN_283; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_285 = 8'h1d == io_inputs_0[7:0] ? 7'h2d : _GEN_284; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_286 = 8'h1e == io_inputs_0[7:0] ? 7'h32 : _GEN_285; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_287 = 8'h1f == io_inputs_0[7:0] ? 7'h37 : _GEN_286; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_288 = 8'h20 == io_inputs_0[7:0] ? 7'h3c : _GEN_287; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_289 = 8'h21 == io_inputs_0[7:0] ? 7'h41 : _GEN_288; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_290 = 8'h22 == io_inputs_0[7:0] ? 7'h46 : _GEN_289; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_291 = 8'h23 == io_inputs_0[7:0] ? 7'h4b : _GEN_290; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_292 = 8'h24 == io_inputs_0[7:0] ? 7'h50 : _GEN_291; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_293 = 8'h25 == io_inputs_0[7:0] ? 7'h55 : _GEN_292; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_294 = 8'h26 == io_inputs_0[7:0] ? 7'h5a : _GEN_293; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_295 = 8'h27 == io_inputs_0[7:0] ? 7'h5f : _GEN_294; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_296 = 8'h28 == io_inputs_0[7:0] ? 7'h64 : _GEN_295; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_297 = 8'h29 == io_inputs_0[7:0] ? 7'h64 : _GEN_296; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_298 = 8'h2a == io_inputs_0[7:0] ? 7'h64 : _GEN_297; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_299 = 8'h2b == io_inputs_0[7:0] ? 7'h64 : _GEN_298; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_300 = 8'h2c == io_inputs_0[7:0] ? 7'h64 : _GEN_299; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_301 = 8'h2d == io_inputs_0[7:0] ? 7'h64 : _GEN_300; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_302 = 8'h2e == io_inputs_0[7:0] ? 7'h64 : _GEN_301; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_303 = 8'h2f == io_inputs_0[7:0] ? 7'h64 : _GEN_302; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_304 = 8'h30 == io_inputs_0[7:0] ? 7'h64 : _GEN_303; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_305 = 8'h31 == io_inputs_0[7:0] ? 7'h64 : _GEN_304; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_306 = 8'h32 == io_inputs_0[7:0] ? 7'h64 : _GEN_305; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_307 = 8'h33 == io_inputs_0[7:0] ? 7'h64 : _GEN_306; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_308 = 8'h34 == io_inputs_0[7:0] ? 7'h64 : _GEN_307; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_309 = 8'h35 == io_inputs_0[7:0] ? 7'h64 : _GEN_308; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_310 = 8'h36 == io_inputs_0[7:0] ? 7'h64 : _GEN_309; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_311 = 8'h37 == io_inputs_0[7:0] ? 7'h64 : _GEN_310; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_312 = 8'h38 == io_inputs_0[7:0] ? 7'h64 : _GEN_311; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_313 = 8'h39 == io_inputs_0[7:0] ? 7'h64 : _GEN_312; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_314 = 8'h3a == io_inputs_0[7:0] ? 7'h64 : _GEN_313; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_315 = 8'h3b == io_inputs_0[7:0] ? 7'h64 : _GEN_314; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_316 = 8'h3c == io_inputs_0[7:0] ? 7'h64 : _GEN_315; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_317 = 8'h3d == io_inputs_0[7:0] ? 7'h5f : _GEN_316; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_318 = 8'h3e == io_inputs_0[7:0] ? 7'h5a : _GEN_317; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_319 = 8'h3f == io_inputs_0[7:0] ? 7'h55 : _GEN_318; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_320 = 8'h40 == io_inputs_0[7:0] ? 7'h50 : _GEN_319; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_321 = 8'h41 == io_inputs_0[7:0] ? 7'h4b : _GEN_320; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_322 = 8'h42 == io_inputs_0[7:0] ? 7'h46 : _GEN_321; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_323 = 8'h43 == io_inputs_0[7:0] ? 7'h41 : _GEN_322; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_324 = 8'h44 == io_inputs_0[7:0] ? 7'h3c : _GEN_323; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_325 = 8'h45 == io_inputs_0[7:0] ? 7'h37 : _GEN_324; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_326 = 8'h46 == io_inputs_0[7:0] ? 7'h32 : _GEN_325; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_327 = 8'h47 == io_inputs_0[7:0] ? 7'h2d : _GEN_326; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_328 = 8'h48 == io_inputs_0[7:0] ? 7'h28 : _GEN_327; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_329 = 8'h49 == io_inputs_0[7:0] ? 7'h23 : _GEN_328; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_330 = 8'h4a == io_inputs_0[7:0] ? 7'h1e : _GEN_329; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_331 = 8'h4b == io_inputs_0[7:0] ? 7'h19 : _GEN_330; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_332 = 8'h4c == io_inputs_0[7:0] ? 7'h14 : _GEN_331; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_333 = 8'h4d == io_inputs_0[7:0] ? 7'hf : _GEN_332; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_334 = 8'h4e == io_inputs_0[7:0] ? 7'ha : _GEN_333; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_335 = 8'h4f == io_inputs_0[7:0] ? 7'h5 : _GEN_334; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_336 = 8'h50 == io_inputs_0[7:0] ? 7'h0 : _GEN_335; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_337 = 8'h51 == io_inputs_0[7:0] ? 7'h0 : _GEN_336; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_338 = 8'h52 == io_inputs_0[7:0] ? 7'h0 : _GEN_337; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_339 = 8'h53 == io_inputs_0[7:0] ? 7'h0 : _GEN_338; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_340 = 8'h54 == io_inputs_0[7:0] ? 7'h0 : _GEN_339; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_341 = 8'h55 == io_inputs_0[7:0] ? 7'h0 : _GEN_340; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_342 = 8'h56 == io_inputs_0[7:0] ? 7'h0 : _GEN_341; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_343 = 8'h57 == io_inputs_0[7:0] ? 7'h0 : _GEN_342; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_344 = 8'h58 == io_inputs_0[7:0] ? 7'h0 : _GEN_343; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_345 = 8'h59 == io_inputs_0[7:0] ? 7'h0 : _GEN_344; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_346 = 8'h5a == io_inputs_0[7:0] ? 7'h0 : _GEN_345; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_347 = 8'h5b == io_inputs_0[7:0] ? 7'h0 : _GEN_346; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_348 = 8'h5c == io_inputs_0[7:0] ? 7'h0 : _GEN_347; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_349 = 8'h5d == io_inputs_0[7:0] ? 7'h0 : _GEN_348; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_350 = 8'h5e == io_inputs_0[7:0] ? 7'h0 : _GEN_349; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_351 = 8'h5f == io_inputs_0[7:0] ? 7'h0 : _GEN_350; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_352 = 8'h60 == io_inputs_0[7:0] ? 7'h0 : _GEN_351; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_353 = 8'h61 == io_inputs_0[7:0] ? 7'h0 : _GEN_352; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_354 = 8'h62 == io_inputs_0[7:0] ? 7'h0 : _GEN_353; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_355 = 8'h63 == io_inputs_0[7:0] ? 7'h0 : _GEN_354; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_356 = 8'h64 == io_inputs_0[7:0] ? 7'h0 : _GEN_355; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_357 = 8'h65 == io_inputs_0[7:0] ? 7'h0 : _GEN_356; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_358 = 8'h66 == io_inputs_0[7:0] ? 7'h0 : _GEN_357; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_359 = 8'h67 == io_inputs_0[7:0] ? 7'h0 : _GEN_358; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_360 = 8'h68 == io_inputs_0[7:0] ? 7'h0 : _GEN_359; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_361 = 8'h69 == io_inputs_0[7:0] ? 7'h0 : _GEN_360; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_362 = 8'h6a == io_inputs_0[7:0] ? 7'h0 : _GEN_361; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_363 = 8'h6b == io_inputs_0[7:0] ? 7'h0 : _GEN_362; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_364 = 8'h6c == io_inputs_0[7:0] ? 7'h0 : _GEN_363; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_365 = 8'h6d == io_inputs_0[7:0] ? 7'h0 : _GEN_364; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_366 = 8'h6e == io_inputs_0[7:0] ? 7'h0 : _GEN_365; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_367 = 8'h6f == io_inputs_0[7:0] ? 7'h0 : _GEN_366; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_368 = 8'h70 == io_inputs_0[7:0] ? 7'h0 : _GEN_367; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_369 = 8'h71 == io_inputs_0[7:0] ? 7'h0 : _GEN_368; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_370 = 8'h72 == io_inputs_0[7:0] ? 7'h0 : _GEN_369; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_371 = 8'h73 == io_inputs_0[7:0] ? 7'h0 : _GEN_370; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_372 = 8'h74 == io_inputs_0[7:0] ? 7'h0 : _GEN_371; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_373 = 8'h75 == io_inputs_0[7:0] ? 7'h0 : _GEN_372; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_374 = 8'h76 == io_inputs_0[7:0] ? 7'h0 : _GEN_373; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_375 = 8'h77 == io_inputs_0[7:0] ? 7'h0 : _GEN_374; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_376 = 8'h78 == io_inputs_0[7:0] ? 7'h0 : _GEN_375; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_377 = 8'h79 == io_inputs_0[7:0] ? 7'h0 : _GEN_376; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_378 = 8'h7a == io_inputs_0[7:0] ? 7'h0 : _GEN_377; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_379 = 8'h7b == io_inputs_0[7:0] ? 7'h0 : _GEN_378; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_380 = 8'h7c == io_inputs_0[7:0] ? 7'h0 : _GEN_379; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_381 = 8'h7d == io_inputs_0[7:0] ? 7'h0 : _GEN_380; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_382 = 8'h7e == io_inputs_0[7:0] ? 7'h0 : _GEN_381; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_383 = 8'h7f == io_inputs_0[7:0] ? 7'h0 : _GEN_382; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_384 = 8'h80 == io_inputs_0[7:0] ? 7'h0 : _GEN_383; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_385 = 8'h81 == io_inputs_0[7:0] ? 7'h0 : _GEN_384; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_386 = 8'h82 == io_inputs_0[7:0] ? 7'h0 : _GEN_385; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_387 = 8'h83 == io_inputs_0[7:0] ? 7'h0 : _GEN_386; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_388 = 8'h84 == io_inputs_0[7:0] ? 7'h0 : _GEN_387; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_389 = 8'h85 == io_inputs_0[7:0] ? 7'h0 : _GEN_388; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_390 = 8'h86 == io_inputs_0[7:0] ? 7'h0 : _GEN_389; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_391 = 8'h87 == io_inputs_0[7:0] ? 7'h0 : _GEN_390; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_392 = 8'h88 == io_inputs_0[7:0] ? 7'h0 : _GEN_391; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_393 = 8'h89 == io_inputs_0[7:0] ? 7'h0 : _GEN_392; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_394 = 8'h8a == io_inputs_0[7:0] ? 7'h0 : _GEN_393; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_395 = 8'h8b == io_inputs_0[7:0] ? 7'h0 : _GEN_394; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_396 = 8'h8c == io_inputs_0[7:0] ? 7'h0 : _GEN_395; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_397 = 8'h8d == io_inputs_0[7:0] ? 7'h0 : _GEN_396; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_398 = 8'h8e == io_inputs_0[7:0] ? 7'h0 : _GEN_397; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_399 = 8'h8f == io_inputs_0[7:0] ? 7'h0 : _GEN_398; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_400 = 8'h90 == io_inputs_0[7:0] ? 7'h0 : _GEN_399; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_401 = 8'h91 == io_inputs_0[7:0] ? 7'h0 : _GEN_400; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_402 = 8'h92 == io_inputs_0[7:0] ? 7'h0 : _GEN_401; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_403 = 8'h93 == io_inputs_0[7:0] ? 7'h0 : _GEN_402; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_404 = 8'h94 == io_inputs_0[7:0] ? 7'h0 : _GEN_403; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_405 = 8'h95 == io_inputs_0[7:0] ? 7'h0 : _GEN_404; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_406 = 8'h96 == io_inputs_0[7:0] ? 7'h0 : _GEN_405; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_407 = 8'h97 == io_inputs_0[7:0] ? 7'h0 : _GEN_406; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_408 = 8'h98 == io_inputs_0[7:0] ? 7'h0 : _GEN_407; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_409 = 8'h99 == io_inputs_0[7:0] ? 7'h0 : _GEN_408; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_410 = 8'h9a == io_inputs_0[7:0] ? 7'h0 : _GEN_409; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_411 = 8'h9b == io_inputs_0[7:0] ? 7'h0 : _GEN_410; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_412 = 8'h9c == io_inputs_0[7:0] ? 7'h0 : _GEN_411; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_413 = 8'h9d == io_inputs_0[7:0] ? 7'h0 : _GEN_412; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_414 = 8'h9e == io_inputs_0[7:0] ? 7'h0 : _GEN_413; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_415 = 8'h9f == io_inputs_0[7:0] ? 7'h0 : _GEN_414; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_416 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_415; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_417 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_416; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_418 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_417; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_419 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_418; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_420 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_419; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_421 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_420; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_422 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_421; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_423 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_422; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_424 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_423; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_425 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_424; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_426 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_425; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_427 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_426; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_428 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_427; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_429 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_428; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_430 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_429; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_431 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_430; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_432 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_431; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_433 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_432; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_434 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_433; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_435 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_434; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_436 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_435; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_437 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_436; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_438 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_437; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_439 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_438; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_440 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_439; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_441 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_440; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_442 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_441; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_443 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_442; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_444 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_443; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_445 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_444; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_446 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_445; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_447 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_446; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_448 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_447; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_449 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_448; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_450 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_449; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_451 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_450; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_452 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_451; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_453 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_452; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_454 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_453; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_455 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_454; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_456 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_455; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_457 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_456; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_458 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_457; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_459 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_458; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_460 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_459; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_461 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_460; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_462 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_461; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_463 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_462; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_464 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_463; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_465 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_464; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_466 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_465; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_467 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_466; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_468 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_467; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_469 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_468; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_470 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_469; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_471 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_470; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_472 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_471; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_473 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_472; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_474 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_473; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_475 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_474; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_476 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_475; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_477 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_476; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_478 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_477; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_479 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_478; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_480 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_479; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_481 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_480; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_482 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_481; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_483 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_482; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_484 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_483; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_485 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_484; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_486 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_485; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_487 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_486; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_488 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_487; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_489 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_488; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_490 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_489; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_491 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_490; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_492 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_491; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_493 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_492; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_494 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_493; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_495 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_494; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_496 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_495; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_497 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_496; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_498 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_497; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_499 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_498; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_500 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_499; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_501 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_500; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_502 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_501; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_503 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_502; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_504 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_503; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_505 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_504; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_506 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_505; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_507 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_506; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_508 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_507; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_509 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_508; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_510 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_509; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_511 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_510; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_573 = 8'h3d == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_574 = 8'h3e == io_inputs_0[7:0] ? 7'ha : _GEN_573; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_575 = 8'h3f == io_inputs_0[7:0] ? 7'hf : _GEN_574; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_576 = 8'h40 == io_inputs_0[7:0] ? 7'h14 : _GEN_575; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_577 = 8'h41 == io_inputs_0[7:0] ? 7'h19 : _GEN_576; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_578 = 8'h42 == io_inputs_0[7:0] ? 7'h1e : _GEN_577; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_579 = 8'h43 == io_inputs_0[7:0] ? 7'h23 : _GEN_578; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_580 = 8'h44 == io_inputs_0[7:0] ? 7'h28 : _GEN_579; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_581 = 8'h45 == io_inputs_0[7:0] ? 7'h2d : _GEN_580; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_582 = 8'h46 == io_inputs_0[7:0] ? 7'h32 : _GEN_581; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_583 = 8'h47 == io_inputs_0[7:0] ? 7'h37 : _GEN_582; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_584 = 8'h48 == io_inputs_0[7:0] ? 7'h3c : _GEN_583; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_585 = 8'h49 == io_inputs_0[7:0] ? 7'h41 : _GEN_584; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_586 = 8'h4a == io_inputs_0[7:0] ? 7'h46 : _GEN_585; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_587 = 8'h4b == io_inputs_0[7:0] ? 7'h4b : _GEN_586; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_588 = 8'h4c == io_inputs_0[7:0] ? 7'h50 : _GEN_587; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_589 = 8'h4d == io_inputs_0[7:0] ? 7'h55 : _GEN_588; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_590 = 8'h4e == io_inputs_0[7:0] ? 7'h5a : _GEN_589; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_591 = 8'h4f == io_inputs_0[7:0] ? 7'h5f : _GEN_590; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_592 = 8'h50 == io_inputs_0[7:0] ? 7'h64 : _GEN_591; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_593 = 8'h51 == io_inputs_0[7:0] ? 7'h64 : _GEN_592; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_594 = 8'h52 == io_inputs_0[7:0] ? 7'h64 : _GEN_593; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_595 = 8'h53 == io_inputs_0[7:0] ? 7'h64 : _GEN_594; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_596 = 8'h54 == io_inputs_0[7:0] ? 7'h64 : _GEN_595; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_597 = 8'h55 == io_inputs_0[7:0] ? 7'h64 : _GEN_596; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_598 = 8'h56 == io_inputs_0[7:0] ? 7'h64 : _GEN_597; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_599 = 8'h57 == io_inputs_0[7:0] ? 7'h64 : _GEN_598; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_600 = 8'h58 == io_inputs_0[7:0] ? 7'h64 : _GEN_599; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_601 = 8'h59 == io_inputs_0[7:0] ? 7'h64 : _GEN_600; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_602 = 8'h5a == io_inputs_0[7:0] ? 7'h64 : _GEN_601; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_603 = 8'h5b == io_inputs_0[7:0] ? 7'h64 : _GEN_602; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_604 = 8'h5c == io_inputs_0[7:0] ? 7'h64 : _GEN_603; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_605 = 8'h5d == io_inputs_0[7:0] ? 7'h64 : _GEN_604; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_606 = 8'h5e == io_inputs_0[7:0] ? 7'h64 : _GEN_605; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_607 = 8'h5f == io_inputs_0[7:0] ? 7'h64 : _GEN_606; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_608 = 8'h60 == io_inputs_0[7:0] ? 7'h64 : _GEN_607; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_609 = 8'h61 == io_inputs_0[7:0] ? 7'h64 : _GEN_608; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_610 = 8'h62 == io_inputs_0[7:0] ? 7'h64 : _GEN_609; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_611 = 8'h63 == io_inputs_0[7:0] ? 7'h64 : _GEN_610; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_612 = 8'h64 == io_inputs_0[7:0] ? 7'h64 : _GEN_611; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_613 = 8'h65 == io_inputs_0[7:0] ? 7'h5f : _GEN_612; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_614 = 8'h66 == io_inputs_0[7:0] ? 7'h5a : _GEN_613; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_615 = 8'h67 == io_inputs_0[7:0] ? 7'h55 : _GEN_614; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_616 = 8'h68 == io_inputs_0[7:0] ? 7'h50 : _GEN_615; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_617 = 8'h69 == io_inputs_0[7:0] ? 7'h4b : _GEN_616; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_618 = 8'h6a == io_inputs_0[7:0] ? 7'h46 : _GEN_617; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_619 = 8'h6b == io_inputs_0[7:0] ? 7'h41 : _GEN_618; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_620 = 8'h6c == io_inputs_0[7:0] ? 7'h3c : _GEN_619; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_621 = 8'h6d == io_inputs_0[7:0] ? 7'h37 : _GEN_620; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_622 = 8'h6e == io_inputs_0[7:0] ? 7'h32 : _GEN_621; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_623 = 8'h6f == io_inputs_0[7:0] ? 7'h2d : _GEN_622; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_624 = 8'h70 == io_inputs_0[7:0] ? 7'h28 : _GEN_623; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_625 = 8'h71 == io_inputs_0[7:0] ? 7'h23 : _GEN_624; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_626 = 8'h72 == io_inputs_0[7:0] ? 7'h1e : _GEN_625; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_627 = 8'h73 == io_inputs_0[7:0] ? 7'h19 : _GEN_626; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_628 = 8'h74 == io_inputs_0[7:0] ? 7'h14 : _GEN_627; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_629 = 8'h75 == io_inputs_0[7:0] ? 7'hf : _GEN_628; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_630 = 8'h76 == io_inputs_0[7:0] ? 7'ha : _GEN_629; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_631 = 8'h77 == io_inputs_0[7:0] ? 7'h5 : _GEN_630; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_632 = 8'h78 == io_inputs_0[7:0] ? 7'h0 : _GEN_631; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_633 = 8'h79 == io_inputs_0[7:0] ? 7'h0 : _GEN_632; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_634 = 8'h7a == io_inputs_0[7:0] ? 7'h0 : _GEN_633; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_635 = 8'h7b == io_inputs_0[7:0] ? 7'h0 : _GEN_634; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_636 = 8'h7c == io_inputs_0[7:0] ? 7'h0 : _GEN_635; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_637 = 8'h7d == io_inputs_0[7:0] ? 7'h0 : _GEN_636; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_638 = 8'h7e == io_inputs_0[7:0] ? 7'h0 : _GEN_637; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_639 = 8'h7f == io_inputs_0[7:0] ? 7'h0 : _GEN_638; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_640 = 8'h80 == io_inputs_0[7:0] ? 7'h0 : _GEN_639; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_641 = 8'h81 == io_inputs_0[7:0] ? 7'h0 : _GEN_640; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_642 = 8'h82 == io_inputs_0[7:0] ? 7'h0 : _GEN_641; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_643 = 8'h83 == io_inputs_0[7:0] ? 7'h0 : _GEN_642; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_644 = 8'h84 == io_inputs_0[7:0] ? 7'h0 : _GEN_643; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_645 = 8'h85 == io_inputs_0[7:0] ? 7'h0 : _GEN_644; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_646 = 8'h86 == io_inputs_0[7:0] ? 7'h0 : _GEN_645; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_647 = 8'h87 == io_inputs_0[7:0] ? 7'h0 : _GEN_646; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_648 = 8'h88 == io_inputs_0[7:0] ? 7'h0 : _GEN_647; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_649 = 8'h89 == io_inputs_0[7:0] ? 7'h0 : _GEN_648; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_650 = 8'h8a == io_inputs_0[7:0] ? 7'h0 : _GEN_649; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_651 = 8'h8b == io_inputs_0[7:0] ? 7'h0 : _GEN_650; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_652 = 8'h8c == io_inputs_0[7:0] ? 7'h0 : _GEN_651; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_653 = 8'h8d == io_inputs_0[7:0] ? 7'h0 : _GEN_652; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_654 = 8'h8e == io_inputs_0[7:0] ? 7'h0 : _GEN_653; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_655 = 8'h8f == io_inputs_0[7:0] ? 7'h0 : _GEN_654; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_656 = 8'h90 == io_inputs_0[7:0] ? 7'h0 : _GEN_655; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_657 = 8'h91 == io_inputs_0[7:0] ? 7'h0 : _GEN_656; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_658 = 8'h92 == io_inputs_0[7:0] ? 7'h0 : _GEN_657; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_659 = 8'h93 == io_inputs_0[7:0] ? 7'h0 : _GEN_658; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_660 = 8'h94 == io_inputs_0[7:0] ? 7'h0 : _GEN_659; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_661 = 8'h95 == io_inputs_0[7:0] ? 7'h0 : _GEN_660; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_662 = 8'h96 == io_inputs_0[7:0] ? 7'h0 : _GEN_661; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_663 = 8'h97 == io_inputs_0[7:0] ? 7'h0 : _GEN_662; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_664 = 8'h98 == io_inputs_0[7:0] ? 7'h0 : _GEN_663; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_665 = 8'h99 == io_inputs_0[7:0] ? 7'h0 : _GEN_664; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_666 = 8'h9a == io_inputs_0[7:0] ? 7'h0 : _GEN_665; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_667 = 8'h9b == io_inputs_0[7:0] ? 7'h0 : _GEN_666; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_668 = 8'h9c == io_inputs_0[7:0] ? 7'h0 : _GEN_667; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_669 = 8'h9d == io_inputs_0[7:0] ? 7'h0 : _GEN_668; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_670 = 8'h9e == io_inputs_0[7:0] ? 7'h0 : _GEN_669; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_671 = 8'h9f == io_inputs_0[7:0] ? 7'h0 : _GEN_670; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_672 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_671; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_673 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_672; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_674 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_673; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_675 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_674; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_676 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_675; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_677 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_676; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_678 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_677; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_679 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_678; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_680 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_679; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_681 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_680; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_682 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_681; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_683 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_682; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_684 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_683; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_685 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_684; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_686 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_685; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_687 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_686; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_688 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_687; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_689 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_688; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_690 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_689; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_691 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_690; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_692 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_691; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_693 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_692; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_694 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_693; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_695 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_694; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_696 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_695; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_697 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_696; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_698 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_697; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_699 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_698; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_700 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_699; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_701 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_700; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_702 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_701; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_703 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_702; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_704 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_703; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_705 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_704; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_706 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_705; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_707 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_706; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_708 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_707; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_709 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_708; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_710 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_709; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_711 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_710; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_712 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_711; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_713 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_712; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_714 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_713; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_715 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_714; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_716 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_715; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_717 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_716; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_718 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_717; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_719 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_718; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_720 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_719; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_721 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_720; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_722 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_721; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_723 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_722; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_724 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_723; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_725 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_724; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_726 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_725; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_727 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_726; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_728 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_727; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_729 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_728; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_730 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_729; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_731 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_730; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_732 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_731; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_733 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_732; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_734 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_733; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_735 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_734; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_736 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_735; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_737 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_736; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_738 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_737; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_739 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_738; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_740 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_739; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_741 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_740; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_742 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_741; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_743 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_742; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_744 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_743; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_745 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_744; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_746 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_745; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_747 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_746; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_748 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_747; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_749 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_748; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_750 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_749; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_751 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_750; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_752 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_751; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_753 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_752; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_754 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_753; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_755 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_754; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_756 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_755; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_757 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_756; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_758 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_757; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_759 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_758; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_760 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_759; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_761 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_760; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_762 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_761; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_763 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_762; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_764 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_763; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_765 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_764; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_766 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_765; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_767 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_766; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_869 = 8'h65 == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_870 = 8'h66 == io_inputs_0[7:0] ? 7'ha : _GEN_869; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_871 = 8'h67 == io_inputs_0[7:0] ? 7'hf : _GEN_870; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_872 = 8'h68 == io_inputs_0[7:0] ? 7'h14 : _GEN_871; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_873 = 8'h69 == io_inputs_0[7:0] ? 7'h19 : _GEN_872; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_874 = 8'h6a == io_inputs_0[7:0] ? 7'h1e : _GEN_873; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_875 = 8'h6b == io_inputs_0[7:0] ? 7'h23 : _GEN_874; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_876 = 8'h6c == io_inputs_0[7:0] ? 7'h28 : _GEN_875; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_877 = 8'h6d == io_inputs_0[7:0] ? 7'h2d : _GEN_876; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_878 = 8'h6e == io_inputs_0[7:0] ? 7'h32 : _GEN_877; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_879 = 8'h6f == io_inputs_0[7:0] ? 7'h37 : _GEN_878; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_880 = 8'h70 == io_inputs_0[7:0] ? 7'h3c : _GEN_879; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_881 = 8'h71 == io_inputs_0[7:0] ? 7'h41 : _GEN_880; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_882 = 8'h72 == io_inputs_0[7:0] ? 7'h46 : _GEN_881; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_883 = 8'h73 == io_inputs_0[7:0] ? 7'h4b : _GEN_882; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_884 = 8'h74 == io_inputs_0[7:0] ? 7'h50 : _GEN_883; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_885 = 8'h75 == io_inputs_0[7:0] ? 7'h55 : _GEN_884; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_886 = 8'h76 == io_inputs_0[7:0] ? 7'h5a : _GEN_885; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_887 = 8'h77 == io_inputs_0[7:0] ? 7'h5f : _GEN_886; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_888 = 8'h78 == io_inputs_0[7:0] ? 7'h64 : _GEN_887; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_889 = 8'h79 == io_inputs_0[7:0] ? 7'h64 : _GEN_888; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_890 = 8'h7a == io_inputs_0[7:0] ? 7'h64 : _GEN_889; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_891 = 8'h7b == io_inputs_0[7:0] ? 7'h64 : _GEN_890; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_892 = 8'h7c == io_inputs_0[7:0] ? 7'h64 : _GEN_891; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_893 = 8'h7d == io_inputs_0[7:0] ? 7'h64 : _GEN_892; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_894 = 8'h7e == io_inputs_0[7:0] ? 7'h64 : _GEN_893; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_895 = 8'h7f == io_inputs_0[7:0] ? 7'h64 : _GEN_894; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_896 = 8'h80 == io_inputs_0[7:0] ? 7'h64 : _GEN_895; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_897 = 8'h81 == io_inputs_0[7:0] ? 7'h64 : _GEN_896; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_898 = 8'h82 == io_inputs_0[7:0] ? 7'h64 : _GEN_897; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_899 = 8'h83 == io_inputs_0[7:0] ? 7'h64 : _GEN_898; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_900 = 8'h84 == io_inputs_0[7:0] ? 7'h64 : _GEN_899; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_901 = 8'h85 == io_inputs_0[7:0] ? 7'h64 : _GEN_900; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_902 = 8'h86 == io_inputs_0[7:0] ? 7'h64 : _GEN_901; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_903 = 8'h87 == io_inputs_0[7:0] ? 7'h64 : _GEN_902; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_904 = 8'h88 == io_inputs_0[7:0] ? 7'h64 : _GEN_903; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_905 = 8'h89 == io_inputs_0[7:0] ? 7'h64 : _GEN_904; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_906 = 8'h8a == io_inputs_0[7:0] ? 7'h64 : _GEN_905; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_907 = 8'h8b == io_inputs_0[7:0] ? 7'h64 : _GEN_906; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_908 = 8'h8c == io_inputs_0[7:0] ? 7'h64 : _GEN_907; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_909 = 8'h8d == io_inputs_0[7:0] ? 7'h5f : _GEN_908; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_910 = 8'h8e == io_inputs_0[7:0] ? 7'h5a : _GEN_909; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_911 = 8'h8f == io_inputs_0[7:0] ? 7'h55 : _GEN_910; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_912 = 8'h90 == io_inputs_0[7:0] ? 7'h50 : _GEN_911; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_913 = 8'h91 == io_inputs_0[7:0] ? 7'h4b : _GEN_912; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_914 = 8'h92 == io_inputs_0[7:0] ? 7'h46 : _GEN_913; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_915 = 8'h93 == io_inputs_0[7:0] ? 7'h41 : _GEN_914; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_916 = 8'h94 == io_inputs_0[7:0] ? 7'h3c : _GEN_915; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_917 = 8'h95 == io_inputs_0[7:0] ? 7'h37 : _GEN_916; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_918 = 8'h96 == io_inputs_0[7:0] ? 7'h32 : _GEN_917; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_919 = 8'h97 == io_inputs_0[7:0] ? 7'h2d : _GEN_918; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_920 = 8'h98 == io_inputs_0[7:0] ? 7'h28 : _GEN_919; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_921 = 8'h99 == io_inputs_0[7:0] ? 7'h23 : _GEN_920; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_922 = 8'h9a == io_inputs_0[7:0] ? 7'h1e : _GEN_921; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_923 = 8'h9b == io_inputs_0[7:0] ? 7'h19 : _GEN_922; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_924 = 8'h9c == io_inputs_0[7:0] ? 7'h14 : _GEN_923; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_925 = 8'h9d == io_inputs_0[7:0] ? 7'hf : _GEN_924; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_926 = 8'h9e == io_inputs_0[7:0] ? 7'ha : _GEN_925; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_927 = 8'h9f == io_inputs_0[7:0] ? 7'h5 : _GEN_926; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_928 = 8'ha0 == io_inputs_0[7:0] ? 7'h0 : _GEN_927; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_929 = 8'ha1 == io_inputs_0[7:0] ? 7'h0 : _GEN_928; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_930 = 8'ha2 == io_inputs_0[7:0] ? 7'h0 : _GEN_929; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_931 = 8'ha3 == io_inputs_0[7:0] ? 7'h0 : _GEN_930; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_932 = 8'ha4 == io_inputs_0[7:0] ? 7'h0 : _GEN_931; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_933 = 8'ha5 == io_inputs_0[7:0] ? 7'h0 : _GEN_932; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_934 = 8'ha6 == io_inputs_0[7:0] ? 7'h0 : _GEN_933; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_935 = 8'ha7 == io_inputs_0[7:0] ? 7'h0 : _GEN_934; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_936 = 8'ha8 == io_inputs_0[7:0] ? 7'h0 : _GEN_935; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_937 = 8'ha9 == io_inputs_0[7:0] ? 7'h0 : _GEN_936; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_938 = 8'haa == io_inputs_0[7:0] ? 7'h0 : _GEN_937; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_939 = 8'hab == io_inputs_0[7:0] ? 7'h0 : _GEN_938; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_940 = 8'hac == io_inputs_0[7:0] ? 7'h0 : _GEN_939; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_941 = 8'had == io_inputs_0[7:0] ? 7'h0 : _GEN_940; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_942 = 8'hae == io_inputs_0[7:0] ? 7'h0 : _GEN_941; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_943 = 8'haf == io_inputs_0[7:0] ? 7'h0 : _GEN_942; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_944 = 8'hb0 == io_inputs_0[7:0] ? 7'h0 : _GEN_943; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_945 = 8'hb1 == io_inputs_0[7:0] ? 7'h0 : _GEN_944; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_946 = 8'hb2 == io_inputs_0[7:0] ? 7'h0 : _GEN_945; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_947 = 8'hb3 == io_inputs_0[7:0] ? 7'h0 : _GEN_946; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_948 = 8'hb4 == io_inputs_0[7:0] ? 7'h0 : _GEN_947; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_949 = 8'hb5 == io_inputs_0[7:0] ? 7'h0 : _GEN_948; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_950 = 8'hb6 == io_inputs_0[7:0] ? 7'h0 : _GEN_949; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_951 = 8'hb7 == io_inputs_0[7:0] ? 7'h0 : _GEN_950; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_952 = 8'hb8 == io_inputs_0[7:0] ? 7'h0 : _GEN_951; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_953 = 8'hb9 == io_inputs_0[7:0] ? 7'h0 : _GEN_952; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_954 = 8'hba == io_inputs_0[7:0] ? 7'h0 : _GEN_953; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_955 = 8'hbb == io_inputs_0[7:0] ? 7'h0 : _GEN_954; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_956 = 8'hbc == io_inputs_0[7:0] ? 7'h0 : _GEN_955; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_957 = 8'hbd == io_inputs_0[7:0] ? 7'h0 : _GEN_956; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_958 = 8'hbe == io_inputs_0[7:0] ? 7'h0 : _GEN_957; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_959 = 8'hbf == io_inputs_0[7:0] ? 7'h0 : _GEN_958; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_960 = 8'hc0 == io_inputs_0[7:0] ? 7'h0 : _GEN_959; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_961 = 8'hc1 == io_inputs_0[7:0] ? 7'h0 : _GEN_960; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_962 = 8'hc2 == io_inputs_0[7:0] ? 7'h0 : _GEN_961; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_963 = 8'hc3 == io_inputs_0[7:0] ? 7'h0 : _GEN_962; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_964 = 8'hc4 == io_inputs_0[7:0] ? 7'h0 : _GEN_963; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_965 = 8'hc5 == io_inputs_0[7:0] ? 7'h0 : _GEN_964; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_966 = 8'hc6 == io_inputs_0[7:0] ? 7'h0 : _GEN_965; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_967 = 8'hc7 == io_inputs_0[7:0] ? 7'h0 : _GEN_966; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_968 = 8'hc8 == io_inputs_0[7:0] ? 7'h0 : _GEN_967; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_969 = 8'hc9 == io_inputs_0[7:0] ? 7'h0 : _GEN_968; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_970 = 8'hca == io_inputs_0[7:0] ? 7'h0 : _GEN_969; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_971 = 8'hcb == io_inputs_0[7:0] ? 7'h0 : _GEN_970; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_972 = 8'hcc == io_inputs_0[7:0] ? 7'h0 : _GEN_971; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_973 = 8'hcd == io_inputs_0[7:0] ? 7'h0 : _GEN_972; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_974 = 8'hce == io_inputs_0[7:0] ? 7'h0 : _GEN_973; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_975 = 8'hcf == io_inputs_0[7:0] ? 7'h0 : _GEN_974; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_976 = 8'hd0 == io_inputs_0[7:0] ? 7'h0 : _GEN_975; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_977 = 8'hd1 == io_inputs_0[7:0] ? 7'h0 : _GEN_976; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_978 = 8'hd2 == io_inputs_0[7:0] ? 7'h0 : _GEN_977; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_979 = 8'hd3 == io_inputs_0[7:0] ? 7'h0 : _GEN_978; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_980 = 8'hd4 == io_inputs_0[7:0] ? 7'h0 : _GEN_979; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_981 = 8'hd5 == io_inputs_0[7:0] ? 7'h0 : _GEN_980; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_982 = 8'hd6 == io_inputs_0[7:0] ? 7'h0 : _GEN_981; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_983 = 8'hd7 == io_inputs_0[7:0] ? 7'h0 : _GEN_982; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_984 = 8'hd8 == io_inputs_0[7:0] ? 7'h0 : _GEN_983; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_985 = 8'hd9 == io_inputs_0[7:0] ? 7'h0 : _GEN_984; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_986 = 8'hda == io_inputs_0[7:0] ? 7'h0 : _GEN_985; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_987 = 8'hdb == io_inputs_0[7:0] ? 7'h0 : _GEN_986; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_988 = 8'hdc == io_inputs_0[7:0] ? 7'h0 : _GEN_987; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_989 = 8'hdd == io_inputs_0[7:0] ? 7'h0 : _GEN_988; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_990 = 8'hde == io_inputs_0[7:0] ? 7'h0 : _GEN_989; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_991 = 8'hdf == io_inputs_0[7:0] ? 7'h0 : _GEN_990; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_992 = 8'he0 == io_inputs_0[7:0] ? 7'h0 : _GEN_991; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_993 = 8'he1 == io_inputs_0[7:0] ? 7'h0 : _GEN_992; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_994 = 8'he2 == io_inputs_0[7:0] ? 7'h0 : _GEN_993; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_995 = 8'he3 == io_inputs_0[7:0] ? 7'h0 : _GEN_994; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_996 = 8'he4 == io_inputs_0[7:0] ? 7'h0 : _GEN_995; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_997 = 8'he5 == io_inputs_0[7:0] ? 7'h0 : _GEN_996; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_998 = 8'he6 == io_inputs_0[7:0] ? 7'h0 : _GEN_997; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_999 = 8'he7 == io_inputs_0[7:0] ? 7'h0 : _GEN_998; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1000 = 8'he8 == io_inputs_0[7:0] ? 7'h0 : _GEN_999; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1001 = 8'he9 == io_inputs_0[7:0] ? 7'h0 : _GEN_1000; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1002 = 8'hea == io_inputs_0[7:0] ? 7'h0 : _GEN_1001; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1003 = 8'heb == io_inputs_0[7:0] ? 7'h0 : _GEN_1002; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1004 = 8'hec == io_inputs_0[7:0] ? 7'h0 : _GEN_1003; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1005 = 8'hed == io_inputs_0[7:0] ? 7'h0 : _GEN_1004; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1006 = 8'hee == io_inputs_0[7:0] ? 7'h0 : _GEN_1005; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1007 = 8'hef == io_inputs_0[7:0] ? 7'h0 : _GEN_1006; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1008 = 8'hf0 == io_inputs_0[7:0] ? 7'h0 : _GEN_1007; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1009 = 8'hf1 == io_inputs_0[7:0] ? 7'h0 : _GEN_1008; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1010 = 8'hf2 == io_inputs_0[7:0] ? 7'h0 : _GEN_1009; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1011 = 8'hf3 == io_inputs_0[7:0] ? 7'h0 : _GEN_1010; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1012 = 8'hf4 == io_inputs_0[7:0] ? 7'h0 : _GEN_1011; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1013 = 8'hf5 == io_inputs_0[7:0] ? 7'h0 : _GEN_1012; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1014 = 8'hf6 == io_inputs_0[7:0] ? 7'h0 : _GEN_1013; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1015 = 8'hf7 == io_inputs_0[7:0] ? 7'h0 : _GEN_1014; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1016 = 8'hf8 == io_inputs_0[7:0] ? 7'h0 : _GEN_1015; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1017 = 8'hf9 == io_inputs_0[7:0] ? 7'h0 : _GEN_1016; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1018 = 8'hfa == io_inputs_0[7:0] ? 7'h0 : _GEN_1017; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1019 = 8'hfb == io_inputs_0[7:0] ? 7'h0 : _GEN_1018; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1020 = 8'hfc == io_inputs_0[7:0] ? 7'h0 : _GEN_1019; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1021 = 8'hfd == io_inputs_0[7:0] ? 7'h0 : _GEN_1020; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1022 = 8'hfe == io_inputs_0[7:0] ? 7'h0 : _GEN_1021; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1023 = 8'hff == io_inputs_0[7:0] ? 7'h0 : _GEN_1022; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1165 = 8'h8d == io_inputs_0[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1166 = 8'h8e == io_inputs_0[7:0] ? 7'ha : _GEN_1165; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1167 = 8'h8f == io_inputs_0[7:0] ? 7'hf : _GEN_1166; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1168 = 8'h90 == io_inputs_0[7:0] ? 7'h14 : _GEN_1167; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1169 = 8'h91 == io_inputs_0[7:0] ? 7'h19 : _GEN_1168; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1170 = 8'h92 == io_inputs_0[7:0] ? 7'h1e : _GEN_1169; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1171 = 8'h93 == io_inputs_0[7:0] ? 7'h23 : _GEN_1170; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1172 = 8'h94 == io_inputs_0[7:0] ? 7'h28 : _GEN_1171; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1173 = 8'h95 == io_inputs_0[7:0] ? 7'h2d : _GEN_1172; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1174 = 8'h96 == io_inputs_0[7:0] ? 7'h32 : _GEN_1173; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1175 = 8'h97 == io_inputs_0[7:0] ? 7'h37 : _GEN_1174; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1176 = 8'h98 == io_inputs_0[7:0] ? 7'h3c : _GEN_1175; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1177 = 8'h99 == io_inputs_0[7:0] ? 7'h41 : _GEN_1176; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1178 = 8'h9a == io_inputs_0[7:0] ? 7'h46 : _GEN_1177; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1179 = 8'h9b == io_inputs_0[7:0] ? 7'h4b : _GEN_1178; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1180 = 8'h9c == io_inputs_0[7:0] ? 7'h50 : _GEN_1179; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1181 = 8'h9d == io_inputs_0[7:0] ? 7'h55 : _GEN_1180; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1182 = 8'h9e == io_inputs_0[7:0] ? 7'h5a : _GEN_1181; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1183 = 8'h9f == io_inputs_0[7:0] ? 7'h5f : _GEN_1182; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1184 = 8'ha0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1183; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1185 = 8'ha1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1184; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1186 = 8'ha2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1185; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1187 = 8'ha3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1186; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1188 = 8'ha4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1187; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1189 = 8'ha5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1188; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1190 = 8'ha6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1189; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1191 = 8'ha7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1190; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1192 = 8'ha8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1191; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1193 = 8'ha9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1192; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1194 = 8'haa == io_inputs_0[7:0] ? 7'h64 : _GEN_1193; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1195 = 8'hab == io_inputs_0[7:0] ? 7'h64 : _GEN_1194; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1196 = 8'hac == io_inputs_0[7:0] ? 7'h64 : _GEN_1195; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1197 = 8'had == io_inputs_0[7:0] ? 7'h64 : _GEN_1196; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1198 = 8'hae == io_inputs_0[7:0] ? 7'h64 : _GEN_1197; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1199 = 8'haf == io_inputs_0[7:0] ? 7'h64 : _GEN_1198; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1200 = 8'hb0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1199; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1201 = 8'hb1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1200; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1202 = 8'hb2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1201; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1203 = 8'hb3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1202; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1204 = 8'hb4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1203; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1205 = 8'hb5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1204; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1206 = 8'hb6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1205; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1207 = 8'hb7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1206; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1208 = 8'hb8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1207; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1209 = 8'hb9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1208; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1210 = 8'hba == io_inputs_0[7:0] ? 7'h64 : _GEN_1209; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1211 = 8'hbb == io_inputs_0[7:0] ? 7'h64 : _GEN_1210; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1212 = 8'hbc == io_inputs_0[7:0] ? 7'h64 : _GEN_1211; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1213 = 8'hbd == io_inputs_0[7:0] ? 7'h64 : _GEN_1212; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1214 = 8'hbe == io_inputs_0[7:0] ? 7'h64 : _GEN_1213; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1215 = 8'hbf == io_inputs_0[7:0] ? 7'h64 : _GEN_1214; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1216 = 8'hc0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1215; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1217 = 8'hc1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1216; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1218 = 8'hc2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1217; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1219 = 8'hc3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1218; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1220 = 8'hc4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1219; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1221 = 8'hc5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1220; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1222 = 8'hc6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1221; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1223 = 8'hc7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1222; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1224 = 8'hc8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1223; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1225 = 8'hc9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1224; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1226 = 8'hca == io_inputs_0[7:0] ? 7'h64 : _GEN_1225; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1227 = 8'hcb == io_inputs_0[7:0] ? 7'h64 : _GEN_1226; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1228 = 8'hcc == io_inputs_0[7:0] ? 7'h64 : _GEN_1227; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1229 = 8'hcd == io_inputs_0[7:0] ? 7'h64 : _GEN_1228; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1230 = 8'hce == io_inputs_0[7:0] ? 7'h64 : _GEN_1229; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1231 = 8'hcf == io_inputs_0[7:0] ? 7'h64 : _GEN_1230; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1232 = 8'hd0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1231; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1233 = 8'hd1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1232; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1234 = 8'hd2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1233; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1235 = 8'hd3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1234; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1236 = 8'hd4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1235; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1237 = 8'hd5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1236; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1238 = 8'hd6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1237; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1239 = 8'hd7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1238; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1240 = 8'hd8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1239; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1241 = 8'hd9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1240; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1242 = 8'hda == io_inputs_0[7:0] ? 7'h64 : _GEN_1241; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1243 = 8'hdb == io_inputs_0[7:0] ? 7'h64 : _GEN_1242; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1244 = 8'hdc == io_inputs_0[7:0] ? 7'h64 : _GEN_1243; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1245 = 8'hdd == io_inputs_0[7:0] ? 7'h64 : _GEN_1244; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1246 = 8'hde == io_inputs_0[7:0] ? 7'h64 : _GEN_1245; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1247 = 8'hdf == io_inputs_0[7:0] ? 7'h64 : _GEN_1246; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1248 = 8'he0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1247; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1249 = 8'he1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1248; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1250 = 8'he2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1249; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1251 = 8'he3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1250; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1252 = 8'he4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1251; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1253 = 8'he5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1252; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1254 = 8'he6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1253; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1255 = 8'he7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1254; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1256 = 8'he8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1255; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1257 = 8'he9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1256; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1258 = 8'hea == io_inputs_0[7:0] ? 7'h64 : _GEN_1257; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1259 = 8'heb == io_inputs_0[7:0] ? 7'h64 : _GEN_1258; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1260 = 8'hec == io_inputs_0[7:0] ? 7'h64 : _GEN_1259; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1261 = 8'hed == io_inputs_0[7:0] ? 7'h64 : _GEN_1260; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1262 = 8'hee == io_inputs_0[7:0] ? 7'h64 : _GEN_1261; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1263 = 8'hef == io_inputs_0[7:0] ? 7'h64 : _GEN_1262; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1264 = 8'hf0 == io_inputs_0[7:0] ? 7'h64 : _GEN_1263; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1265 = 8'hf1 == io_inputs_0[7:0] ? 7'h64 : _GEN_1264; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1266 = 8'hf2 == io_inputs_0[7:0] ? 7'h64 : _GEN_1265; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1267 = 8'hf3 == io_inputs_0[7:0] ? 7'h64 : _GEN_1266; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1268 = 8'hf4 == io_inputs_0[7:0] ? 7'h64 : _GEN_1267; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1269 = 8'hf5 == io_inputs_0[7:0] ? 7'h64 : _GEN_1268; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1270 = 8'hf6 == io_inputs_0[7:0] ? 7'h64 : _GEN_1269; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1271 = 8'hf7 == io_inputs_0[7:0] ? 7'h64 : _GEN_1270; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1272 = 8'hf8 == io_inputs_0[7:0] ? 7'h64 : _GEN_1271; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1273 = 8'hf9 == io_inputs_0[7:0] ? 7'h64 : _GEN_1272; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1274 = 8'hfa == io_inputs_0[7:0] ? 7'h64 : _GEN_1273; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1275 = 8'hfb == io_inputs_0[7:0] ? 7'h64 : _GEN_1274; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1276 = 8'hfc == io_inputs_0[7:0] ? 7'h64 : _GEN_1275; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1277 = 8'hfd == io_inputs_0[7:0] ? 7'h64 : _GEN_1276; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1278 = 8'hfe == io_inputs_0[7:0] ? 7'h64 : _GEN_1277; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_1279 = 8'hff == io_inputs_0[7:0] ? 7'h64 : _GEN_1278; // @[regular_fuzzification.scala 176:{36,36}]
  wire [6:0] _GEN_6425 = io_start ? _GEN_255 : {{4'd0}, regLutResultsVec_0}; // @[regular_fuzzification.scala 125:29 163:29 176:36]
  wire [6:0] _GEN_6426 = io_start ? _GEN_511 : {{4'd0}, regLutResultsVec_1}; // @[regular_fuzzification.scala 125:29 163:29 176:36]
  wire [6:0] _GEN_6427 = io_start ? _GEN_767 : {{4'd0}, regLutResultsVec_2}; // @[regular_fuzzification.scala 125:29 163:29 176:36]
  wire [6:0] _GEN_6428 = io_start ? _GEN_1023 : {{4'd0}, regLutResultsVec_3}; // @[regular_fuzzification.scala 125:29 163:29 176:36]
  wire [6:0] _GEN_6429 = io_start ? _GEN_1279 : {{4'd0}, regLutResultsVec_4}; // @[regular_fuzzification.scala 125:29 163:29 176:36]
  wire [2:0] regMaxVec_0_result = regMaxVec_0_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_1_result = regMaxVec_1_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_2_result = regMaxVec_2_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_3_result = regMaxVec_3_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] regMaxVec_4_result = regMaxVec_4_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [2:0] outResult_result = outResult_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  MultipleComparator regMaxVec_0_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_0_comparatorModule_clock),
    .io_start(regMaxVec_0_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_0_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_0_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_0_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_0_comparatorModule_io_inputs_3),
    .io_result(regMaxVec_0_comparatorModule_io_result)
  );
  MultipleComparator_1 regMaxVec_1_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_1_comparatorModule_clock),
    .io_start(regMaxVec_1_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_1_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_1_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_1_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_1_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_1_comparatorModule_io_inputs_4),
    .io_inputs_5(regMaxVec_1_comparatorModule_io_inputs_5),
    .io_result(regMaxVec_1_comparatorModule_io_result)
  );
  MultipleComparator regMaxVec_2_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_2_comparatorModule_clock),
    .io_start(regMaxVec_2_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_2_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_2_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_2_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_2_comparatorModule_io_inputs_3),
    .io_result(regMaxVec_2_comparatorModule_io_result)
  );
  MultipleComparator_1 regMaxVec_3_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_3_comparatorModule_clock),
    .io_start(regMaxVec_3_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_3_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_3_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_3_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_3_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_3_comparatorModule_io_inputs_4),
    .io_inputs_5(regMaxVec_3_comparatorModule_io_inputs_5),
    .io_result(regMaxVec_3_comparatorModule_io_result)
  );
  MultipleComparator_4 regMaxVec_4_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_4_comparatorModule_clock),
    .io_start(regMaxVec_4_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_4_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_4_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_4_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_4_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_4_comparatorModule_io_inputs_4),
    .io_result(regMaxVec_4_comparatorModule_io_result)
  );
  MultipleComparator_5 outResult_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(outResult_comparatorModule_clock),
    .io_start(outResult_comparatorModule_io_start),
    .io_inputs_0(outResult_comparatorModule_io_inputs_0),
    .io_inputs_1(outResult_comparatorModule_io_inputs_1),
    .io_inputs_2(outResult_comparatorModule_io_inputs_2),
    .io_inputs_3(outResult_comparatorModule_io_inputs_3),
    .io_inputs_4(outResult_comparatorModule_io_inputs_4),
    .io_result(outResult_comparatorModule_io_result)
  );
  assign io_outResultValid = 1'h0; // @[regular_fuzzification.scala 163:29 404:20]
  assign io_outResult = io_start ? outResult_result : 3'h0; // @[regular_fuzzification.scala 163:29 378:15 403:15]
  assign regMaxVec_0_comparatorModule_clock = clock;
  assign regMaxVec_0_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_0_comparatorModule_io_inputs_0 = regMinVec_0; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_0_comparatorModule_io_inputs_1 = regMinVec_1; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_0_comparatorModule_io_inputs_2 = regMinVec_2; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_0_comparatorModule_io_inputs_3 = regMinVec_5; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_1_comparatorModule_clock = clock;
  assign regMaxVec_1_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_1_comparatorModule_io_inputs_0 = regMinVec_3; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_1_comparatorModule_io_inputs_1 = regMinVec_4; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_1_comparatorModule_io_inputs_2 = regMinVec_6; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_1_comparatorModule_io_inputs_3 = regMinVec_7; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_1_comparatorModule_io_inputs_4 = regMinVec_8; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_1_comparatorModule_io_inputs_5 = regMinVec_10; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_2_comparatorModule_clock = clock;
  assign regMaxVec_2_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_2_comparatorModule_io_inputs_0 = regMinVec_9; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_2_comparatorModule_io_inputs_1 = regMinVec_11; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_2_comparatorModule_io_inputs_2 = regMinVec_12; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_2_comparatorModule_io_inputs_3 = regMinVec_15; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_3_comparatorModule_clock = clock;
  assign regMaxVec_3_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_3_comparatorModule_io_inputs_0 = regMinVec_13; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_3_comparatorModule_io_inputs_1 = regMinVec_14; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_3_comparatorModule_io_inputs_2 = regMinVec_16; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_3_comparatorModule_io_inputs_3 = regMinVec_17; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_3_comparatorModule_io_inputs_4 = regMinVec_20; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_3_comparatorModule_io_inputs_5 = regMinVec_21; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_4_comparatorModule_clock = clock;
  assign regMaxVec_4_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_4_comparatorModule_io_inputs_0 = regMinVec_18; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_4_comparatorModule_io_inputs_1 = regMinVec_19; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_4_comparatorModule_io_inputs_2 = regMinVec_22; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_4_comparatorModule_io_inputs_3 = regMinVec_23; // @[regular_fuzzification.scala 309:15 312:30]
  assign regMaxVec_4_comparatorModule_io_inputs_4 = regMinVec_24; // @[regular_fuzzification.scala 309:15 312:30]
  assign outResult_comparatorModule_clock = clock;
  assign outResult_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign outResult_comparatorModule_io_inputs_0 = regMaxVec_0; // @[regular_fuzzification.scala 361:11 368:40]
  assign outResult_comparatorModule_io_inputs_1 = regMaxVec_1; // @[regular_fuzzification.scala 361:11 368:40]
  assign outResult_comparatorModule_io_inputs_2 = regMaxVec_2; // @[regular_fuzzification.scala 361:11 368:40]
  assign outResult_comparatorModule_io_inputs_3 = regMaxVec_3; // @[regular_fuzzification.scala 361:11 368:40]
  assign outResult_comparatorModule_io_inputs_4 = regMaxVec_4; // @[regular_fuzzification.scala 361:11 368:40]
  always @(posedge clock) begin
    regLutResultsVec_0 <= _GEN_6425[2:0];
    regLutResultsVec_1 <= _GEN_6426[2:0];
    regLutResultsVec_2 <= _GEN_6427[2:0];
    regLutResultsVec_3 <= _GEN_6428[2:0];
    regLutResultsVec_4 <= _GEN_6429[2:0];
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_0 <= regLutResultsVec_0; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_1 <= regLutResultsVec_0; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_2 <= regLutResultsVec_0; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_3 <= regLutResultsVec_0; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_4 <= regLutResultsVec_0; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_5 <= regLutResultsVec_1; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_6 <= regLutResultsVec_1; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_7 <= regLutResultsVec_1; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_8 <= regLutResultsVec_1; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_9 <= regLutResultsVec_1; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_10 <= regLutResultsVec_2; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_11 <= regLutResultsVec_2; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_12 <= regLutResultsVec_2; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_13 <= regLutResultsVec_2; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_14 <= regLutResultsVec_2; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_15 <= regLutResultsVec_3; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_16 <= regLutResultsVec_3; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_17 <= regLutResultsVec_3; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_18 <= regLutResultsVec_3; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_19 <= regLutResultsVec_3; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_20 <= regLutResultsVec_4; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_21 <= regLutResultsVec_4; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_22 <= regLutResultsVec_4; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_23 <= regLutResultsVec_4; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMinVec_24 <= regLutResultsVec_4; // @[regular_fuzzification.scala 247:38]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMaxVec_0 <= regMaxVec_0_result; // @[regular_fuzzification.scala 315:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMaxVec_1 <= regMaxVec_1_result; // @[regular_fuzzification.scala 315:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMaxVec_2 <= regMaxVec_2_result; // @[regular_fuzzification.scala 315:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMaxVec_3 <= regMaxVec_3_result; // @[regular_fuzzification.scala 315:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 163:29]
      regMaxVec_4 <= regMaxVec_4_result; // @[regular_fuzzification.scala 315:39]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_0,regLutResultsVec_0); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_0,regLutResultsVec_0); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_0,regLutResultsVec_0); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_0,regLutResultsVec_0); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_0,regLutResultsVec_0); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_1,regLutResultsVec_1); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_1,regLutResultsVec_1); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_1,regLutResultsVec_1); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_1,regLutResultsVec_1); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_1,regLutResultsVec_1); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_2,regLutResultsVec_2); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_2,regLutResultsVec_2); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_2,regLutResultsVec_2); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_2,regLutResultsVec_2); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_2,regLutResultsVec_2); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_3,regLutResultsVec_3); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_3,regLutResultsVec_3); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_3,regLutResultsVec_3); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_3,regLutResultsVec_3); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_3,regLutResultsVec_3); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_4,regLutResultsVec_4); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_4,regLutResultsVec_4); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_4,regLutResultsVec_4); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_4,regLutResultsVec_4); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_start & ~reset) begin
          $fwrite(32'h80000002,"dbg, regular comparator without index | start : %d | input1 : %d, input2 : %d\n",
            io_start,regLutResultsVec_4,regLutResultsVec_4); // @[comparator.scala 82:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
