module Comparator(
  input  [6:0] io_in1,
  input  [6:0] io_in2,
  output       io_maxMin
);
  assign io_maxMin = io_in1 >= io_in2; // @[comparator.scala 34:15]
endmodule
module Comparator_25(
  input  [6:0] io_in1,
  input  [6:0] io_in2,
  output       io_maxMin
);
  assign io_maxMin = io_in1 >= io_in2 ? 1'h0 : 1'h1; // @[comparator.scala 34:26 37:20 45:20]
endmodule
module MultipleComparator(
  input        clock,
  input        io_start,
  input  [6:0] io_inputs_0,
  input  [6:0] io_inputs_1,
  input  [6:0] io_inputs_2,
  input  [6:0] io_inputs_3,
  output [6:0] io_result
);
  wire [6:0] regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  reg [6:0] regMinMaxResultVec_0_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_1_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_2_minMaxResult; // @[multiple_comparator.scala 113:31]
  wire  regMinMaxResultVec_0_minMaxResult_maxMinOutput = regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_1_minMaxResult_maxMinOutput = regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_2_minMaxResult_maxMinOutput = regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  Comparator_25 regMinMaxResultVec_0_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_1_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_2_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin)
  );
  assign io_result = regMinMaxResultVec_2_minMaxResult; // @[multiple_comparator.scala 274:13]
  assign regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1 = io_inputs_0; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2 = io_inputs_1; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1 = io_inputs_2; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2 = io_inputs_3; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1 = regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2 = regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 77:29]
  always @(posedge clock) begin
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_0_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_0_minMaxResult <= io_inputs_0; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_0_minMaxResult <= io_inputs_1; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_1_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_1_minMaxResult <= io_inputs_2; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_1_minMaxResult <= io_inputs_3; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_2_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_2_minMaxResult <= regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_2_minMaxResult <= regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 103:14]
      end
    end
  end
endmodule
module MultipleComparator_1(
  input        clock,
  input        io_start,
  input  [6:0] io_inputs_0,
  input  [6:0] io_inputs_1,
  input  [6:0] io_inputs_2,
  input  [6:0] io_inputs_3,
  input  [6:0] io_inputs_4,
  input  [6:0] io_inputs_5,
  output [6:0] io_result
);
  wire [6:0] regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_3_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_4_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_4_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_4_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  reg [6:0] regMinMaxResultVec_0_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_1_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_2_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_3_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_4_minMaxResult; // @[multiple_comparator.scala 113:31]
  wire  regMinMaxResultVec_0_minMaxResult_maxMinOutput = regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_1_minMaxResult_maxMinOutput = regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_2_minMaxResult_maxMinOutput = regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_3_minMaxResult_maxMinOutput = regMinMaxResultVec_3_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_4_minMaxResult_maxMinOutput = regMinMaxResultVec_4_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  Comparator_25 regMinMaxResultVec_0_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_1_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_2_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_3_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_3_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_4_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_4_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_4_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_4_minMaxResult_comparatorModule_io_maxMin)
  );
  assign io_result = regMinMaxResultVec_4_minMaxResult; // @[multiple_comparator.scala 274:13]
  assign regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1 = io_inputs_0; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2 = io_inputs_1; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1 = io_inputs_2; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2 = io_inputs_3; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1 = io_inputs_4; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2 = io_inputs_5; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in1 = regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in2 = regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_4_minMaxResult_comparatorModule_io_in1 = regMinMaxResultVec_2_minMaxResult; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_4_minMaxResult_comparatorModule_io_in2 = regMinMaxResultVec_3_minMaxResult; // @[comparator.scala 77:29]
  always @(posedge clock) begin
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_0_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_0_minMaxResult <= io_inputs_0; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_0_minMaxResult <= io_inputs_1; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_1_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_1_minMaxResult <= io_inputs_2; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_1_minMaxResult <= io_inputs_3; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_2_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_2_minMaxResult <= io_inputs_4; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_2_minMaxResult <= io_inputs_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_3_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_3_minMaxResult <= regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_3_minMaxResult <= regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_4_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_4_minMaxResult <= regMinMaxResultVec_2_minMaxResult; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_4_minMaxResult <= regMinMaxResultVec_3_minMaxResult; // @[comparator.scala 103:14]
      end
    end
  end
endmodule
module MultipleComparator_4(
  input        clock,
  input        io_start,
  input  [6:0] io_inputs_0,
  input  [6:0] io_inputs_1,
  input  [6:0] io_inputs_2,
  input  [6:0] io_inputs_3,
  input  [6:0] io_inputs_4,
  output [6:0] io_result
);
  wire [6:0] regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinMaxResultVec_3_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  reg [6:0] regMinMaxResultVec_0_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_1_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_2_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_3_minMaxResult; // @[multiple_comparator.scala 113:31]
  wire  regMinMaxResultVec_0_minMaxResult_maxMinOutput = regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_1_minMaxResult_maxMinOutput = regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_2_minMaxResult_maxMinOutput = regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinMaxResultVec_3_minMaxResult_maxMinOutput = regMinMaxResultVec_3_minMaxResult_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  Comparator_25 regMinMaxResultVec_0_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_0_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_1_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_1_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_2_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_2_minMaxResult_comparatorModule_io_maxMin)
  );
  Comparator_25 regMinMaxResultVec_3_minMaxResult_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in1),
    .io_in2(regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in2),
    .io_maxMin(regMinMaxResultVec_3_minMaxResult_comparatorModule_io_maxMin)
  );
  assign io_result = regMinMaxResultVec_3_minMaxResult; // @[multiple_comparator.scala 274:13]
  assign regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in1 = io_inputs_0; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_0_minMaxResult_comparatorModule_io_in2 = io_inputs_1; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in1 = io_inputs_2; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_1_minMaxResult_comparatorModule_io_in2 = io_inputs_3; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in1 = regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_2_minMaxResult_comparatorModule_io_in2 = regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 77:29]
  assign regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in1 = regMinMaxResultVec_2_minMaxResult; // @[comparator.scala 76:29]
  assign regMinMaxResultVec_3_minMaxResult_comparatorModule_io_in2 = io_inputs_4; // @[comparator.scala 77:29]
  always @(posedge clock) begin
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_0_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_0_minMaxResult <= io_inputs_0; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_0_minMaxResult <= io_inputs_1; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_1_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_1_minMaxResult <= io_inputs_2; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_1_minMaxResult <= io_inputs_3; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_2_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_2_minMaxResult <= regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_2_minMaxResult <= regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~regMinMaxResultVec_3_minMaxResult_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinMaxResultVec_3_minMaxResult <= regMinMaxResultVec_2_minMaxResult; // @[comparator.scala 101:14]
      end else begin
        regMinMaxResultVec_3_minMaxResult <= io_inputs_4; // @[comparator.scala 103:14]
      end
    end
  end
endmodule
module MultipleComparator_5(
  input        clock,
  input        io_start,
  input  [6:0] io_inputs_0,
  input  [6:0] io_inputs_1,
  input  [6:0] io_inputs_2,
  input  [6:0] io_inputs_3,
  input  [6:0] io_inputs_4,
  output [6:0] io_result
);
  wire [6:0] comparatorModule_io_in1; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_io_in2; // @[comparator.scala 121:34]
  wire  comparatorModule_io_maxMin; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_1_io_in1; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_1_io_in2; // @[comparator.scala 121:34]
  wire  comparatorModule_1_io_maxMin; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_2_io_in1; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_2_io_in2; // @[comparator.scala 121:34]
  wire  comparatorModule_2_io_maxMin; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_3_io_in1; // @[comparator.scala 121:34]
  wire [6:0] comparatorModule_3_io_in2; // @[comparator.scala 121:34]
  wire  comparatorModule_3_io_maxMin; // @[comparator.scala 121:34]
  reg [6:0] regMinMaxResultVec_0_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [2:0] regMinMaxResultVec_0_minMaxIndex; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_1_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [2:0] regMinMaxResultVec_1_minMaxIndex; // @[multiple_comparator.scala 113:31]
  reg [6:0] regMinMaxResultVec_2_minMaxResult; // @[multiple_comparator.scala 113:31]
  reg [2:0] regMinMaxResultVec_2_minMaxIndex; // @[multiple_comparator.scala 113:31]
  reg [2:0] regMinMaxResultVec_3_minMaxIndex; // @[multiple_comparator.scala 113:31]
  wire  maxMinOutput_1 = comparatorModule_io_maxMin; // @[comparator.scala 126:28 145:18]
  wire  _GEN_1 = ~maxMinOutput_1 ? 1'h0 : 1'h1; // @[comparator.scala 155:40 157:19 160:19]
  wire  maxMinOutput_2 = comparatorModule_1_io_maxMin; // @[comparator.scala 126:28 145:18]
  wire [1:0] _GEN_3 = ~maxMinOutput_2 ? 2'h2 : 2'h3; // @[comparator.scala 155:40 157:19 160:19]
  wire  maxMinOutput_3 = comparatorModule_2_io_maxMin; // @[comparator.scala 126:28 145:18]
  wire [2:0] _GEN_5 = ~maxMinOutput_3 ? regMinMaxResultVec_0_minMaxIndex : regMinMaxResultVec_1_minMaxIndex; // @[comparator.scala 155:40 157:19 160:19]
  wire  maxMinOutput_4 = comparatorModule_3_io_maxMin; // @[comparator.scala 126:28 145:18]
  wire [2:0] _GEN_7 = ~maxMinOutput_4 ? regMinMaxResultVec_2_minMaxIndex : 3'h4; // @[comparator.scala 155:40 157:19 160:19]
  wire [6:0] resultIndex = {{6'd0}, _GEN_1}; // @[comparator.scala 124:27]
  wire [6:0] _GEN_9 = io_start ? resultIndex : {{4'd0}, regMinMaxResultVec_0_minMaxIndex}; // @[multiple_comparator.scala 130:18 113:31 170:45]
  wire [6:0] resultIndex_1 = {{5'd0}, _GEN_3}; // @[comparator.scala 124:27]
  wire [6:0] _GEN_11 = io_start ? resultIndex_1 : {{4'd0}, regMinMaxResultVec_1_minMaxIndex}; // @[multiple_comparator.scala 130:18 113:31 170:45]
  wire [6:0] resultIndex_2 = {{4'd0}, _GEN_5}; // @[comparator.scala 124:27]
  wire [6:0] _GEN_13 = io_start ? resultIndex_2 : {{4'd0}, regMinMaxResultVec_2_minMaxIndex}; // @[multiple_comparator.scala 130:18 113:31 249:47]
  wire [6:0] resultIndex_3 = {{4'd0}, _GEN_7}; // @[comparator.scala 124:27]
  wire [6:0] _GEN_15 = io_start ? resultIndex_3 : {{4'd0}, regMinMaxResultVec_3_minMaxIndex}; // @[multiple_comparator.scala 130:18 113:31 214:51]
  Comparator_25 comparatorModule ( // @[comparator.scala 121:34]
    .io_in1(comparatorModule_io_in1),
    .io_in2(comparatorModule_io_in2),
    .io_maxMin(comparatorModule_io_maxMin)
  );
  Comparator_25 comparatorModule_1 ( // @[comparator.scala 121:34]
    .io_in1(comparatorModule_1_io_in1),
    .io_in2(comparatorModule_1_io_in2),
    .io_maxMin(comparatorModule_1_io_maxMin)
  );
  Comparator_25 comparatorModule_2 ( // @[comparator.scala 121:34]
    .io_in1(comparatorModule_2_io_in1),
    .io_in2(comparatorModule_2_io_in2),
    .io_maxMin(comparatorModule_2_io_maxMin)
  );
  Comparator_25 comparatorModule_3 ( // @[comparator.scala 121:34]
    .io_in1(comparatorModule_3_io_in1),
    .io_in2(comparatorModule_3_io_in2),
    .io_maxMin(comparatorModule_3_io_maxMin)
  );
  assign io_result = {{4'd0}, regMinMaxResultVec_3_minMaxIndex}; // @[multiple_comparator.scala 274:13]
  assign comparatorModule_io_in1 = io_inputs_0; // @[comparator.scala 131:29]
  assign comparatorModule_io_in2 = io_inputs_1; // @[comparator.scala 132:29]
  assign comparatorModule_1_io_in1 = io_inputs_2; // @[comparator.scala 131:29]
  assign comparatorModule_1_io_in2 = io_inputs_3; // @[comparator.scala 132:29]
  assign comparatorModule_2_io_in1 = regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 131:29]
  assign comparatorModule_2_io_in2 = regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 132:29]
  assign comparatorModule_3_io_in1 = regMinMaxResultVec_2_minMaxResult; // @[comparator.scala 131:29]
  assign comparatorModule_3_io_in2 = io_inputs_4; // @[comparator.scala 132:29]
  always @(posedge clock) begin
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~maxMinOutput_1) begin // @[comparator.scala 155:40]
        regMinMaxResultVec_0_minMaxResult <= io_inputs_0; // @[comparator.scala 156:14]
      end else begin
        regMinMaxResultVec_0_minMaxResult <= io_inputs_1; // @[comparator.scala 159:14]
      end
    end
    regMinMaxResultVec_0_minMaxIndex <= _GEN_9[2:0];
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~maxMinOutput_2) begin // @[comparator.scala 155:40]
        regMinMaxResultVec_1_minMaxResult <= io_inputs_2; // @[comparator.scala 156:14]
      end else begin
        regMinMaxResultVec_1_minMaxResult <= io_inputs_3; // @[comparator.scala 159:14]
      end
    end
    regMinMaxResultVec_1_minMaxIndex <= _GEN_11[2:0];
    if (io_start) begin // @[multiple_comparator.scala 130:18]
      if (~maxMinOutput_3) begin // @[comparator.scala 155:40]
        regMinMaxResultVec_2_minMaxResult <= regMinMaxResultVec_0_minMaxResult; // @[comparator.scala 156:14]
      end else begin
        regMinMaxResultVec_2_minMaxResult <= regMinMaxResultVec_1_minMaxResult; // @[comparator.scala 159:14]
      end
    end
    regMinMaxResultVec_2_minMaxIndex <= _GEN_13[2:0];
    regMinMaxResultVec_3_minMaxIndex <= _GEN_15[2:0];
  end
endmodule
module RegularFuzzification(
  input        clock,
  input        reset,
  input        io_start,
  input  [9:0] io_inputs_0,
  input  [9:0] io_inputs_1,
  input  [6:0] io_lutConnections_0,
  input  [6:0] io_lutConnections_1,
  input  [6:0] io_lutConnections_2,
  input  [6:0] io_lutConnections_3,
  input  [6:0] io_lutConnections_4,
  input  [6:0] io_lutConnections_5,
  input  [6:0] io_lutConnections_6,
  input  [6:0] io_lutConnections_7,
  input  [6:0] io_lutConnections_8,
  input  [6:0] io_lutConnections_9,
  output       io_outResultValid,
  output [6:0] io_outResult
);
  wire [6:0] regMinVec_0_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_0_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_0_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_1_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_1_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_1_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_2_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_2_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_2_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_3_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_3_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_3_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_4_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_4_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_4_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_5_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_5_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_5_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_6_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_6_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_6_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_7_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_7_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_7_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_8_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_8_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_8_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_9_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_9_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_9_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_10_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_10_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_10_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_11_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_11_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_11_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_12_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_12_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_12_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_13_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_13_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_13_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_14_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_14_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_14_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_15_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_15_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_15_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_16_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_16_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_16_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_17_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_17_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_17_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_18_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_18_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_18_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_19_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_19_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_19_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_20_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_20_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_20_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_21_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_21_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_21_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_22_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_22_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_22_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_23_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_23_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_23_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_24_comparatorModule_io_in1; // @[comparator.scala 69:34]
  wire [6:0] regMinVec_24_comparatorModule_io_in2; // @[comparator.scala 69:34]
  wire  regMinVec_24_comparatorModule_io_maxMin; // @[comparator.scala 69:34]
  wire  regMaxVec_0_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_0_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_0_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_0_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_0_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_0_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_0_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_1_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_1_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_inputs_5; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_1_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_2_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_2_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_2_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_2_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_2_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_2_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_2_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_3_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_3_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_inputs_5; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_3_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_4_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  regMaxVec_4_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_4_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_4_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_4_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_4_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_4_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [6:0] regMaxVec_4_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  wire  outResult_comparatorModule_clock; // @[multiple_comparator.scala 293:34]
  wire  outResult_comparatorModule_io_start; // @[multiple_comparator.scala 293:34]
  wire [6:0] outResult_comparatorModule_io_inputs_0; // @[multiple_comparator.scala 293:34]
  wire [6:0] outResult_comparatorModule_io_inputs_1; // @[multiple_comparator.scala 293:34]
  wire [6:0] outResult_comparatorModule_io_inputs_2; // @[multiple_comparator.scala 293:34]
  wire [6:0] outResult_comparatorModule_io_inputs_3; // @[multiple_comparator.scala 293:34]
  wire [6:0] outResult_comparatorModule_io_inputs_4; // @[multiple_comparator.scala 293:34]
  wire [6:0] outResult_comparatorModule_io_result; // @[multiple_comparator.scala 293:34]
  reg [6:0] regLutResultsVec_0; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_1; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_2; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_3; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_4; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_5; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_6; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_7; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_8; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regLutResultsVec_9; // @[regular_fuzzification.scala 132:29]
  reg [6:0] regMinVec_0; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_1; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_2; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_3; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_4; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_5; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_6; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_7; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_8; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_9; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_10; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_11; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_12; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_13; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_14; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_15; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_16; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_17; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_18; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_19; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_20; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_21; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_22; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_23; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMinVec_24; // @[regular_fuzzification.scala 151:22]
  reg [6:0] regMaxVec_0; // @[regular_fuzzification.scala 166:22]
  reg [6:0] regMaxVec_1; // @[regular_fuzzification.scala 166:22]
  reg [6:0] regMaxVec_2; // @[regular_fuzzification.scala 166:22]
  reg [6:0] regMaxVec_3; // @[regular_fuzzification.scala 166:22]
  reg [6:0] regMaxVec_4; // @[regular_fuzzification.scala 166:22]
  wire [6:0] _GEN_51 = 10'h33 == io_inputs_0 ? 7'h63 : 7'h64; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_52 = 10'h34 == io_inputs_0 ? 7'h62 : _GEN_51; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_53 = 10'h35 == io_inputs_0 ? 7'h61 : _GEN_52; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_54 = 10'h36 == io_inputs_0 ? 7'h60 : _GEN_53; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_55 = 10'h37 == io_inputs_0 ? 7'h5f : _GEN_54; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_56 = 10'h38 == io_inputs_0 ? 7'h5e : _GEN_55; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_57 = 10'h39 == io_inputs_0 ? 7'h5d : _GEN_56; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_58 = 10'h3a == io_inputs_0 ? 7'h5c : _GEN_57; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_59 = 10'h3b == io_inputs_0 ? 7'h5b : _GEN_58; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_60 = 10'h3c == io_inputs_0 ? 7'h5a : _GEN_59; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_61 = 10'h3d == io_inputs_0 ? 7'h59 : _GEN_60; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_62 = 10'h3e == io_inputs_0 ? 7'h58 : _GEN_61; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_63 = 10'h3f == io_inputs_0 ? 7'h57 : _GEN_62; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_64 = 10'h40 == io_inputs_0 ? 7'h56 : _GEN_63; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_65 = 10'h41 == io_inputs_0 ? 7'h55 : _GEN_64; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_66 = 10'h42 == io_inputs_0 ? 7'h54 : _GEN_65; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_67 = 10'h43 == io_inputs_0 ? 7'h53 : _GEN_66; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_68 = 10'h44 == io_inputs_0 ? 7'h52 : _GEN_67; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_69 = 10'h45 == io_inputs_0 ? 7'h51 : _GEN_68; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_70 = 10'h46 == io_inputs_0 ? 7'h50 : _GEN_69; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_71 = 10'h47 == io_inputs_0 ? 7'h4f : _GEN_70; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_72 = 10'h48 == io_inputs_0 ? 7'h4e : _GEN_71; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_73 = 10'h49 == io_inputs_0 ? 7'h4d : _GEN_72; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_74 = 10'h4a == io_inputs_0 ? 7'h4c : _GEN_73; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_75 = 10'h4b == io_inputs_0 ? 7'h4b : _GEN_74; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_76 = 10'h4c == io_inputs_0 ? 7'h4a : _GEN_75; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_77 = 10'h4d == io_inputs_0 ? 7'h49 : _GEN_76; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_78 = 10'h4e == io_inputs_0 ? 7'h48 : _GEN_77; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_79 = 10'h4f == io_inputs_0 ? 7'h47 : _GEN_78; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_80 = 10'h50 == io_inputs_0 ? 7'h46 : _GEN_79; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_81 = 10'h51 == io_inputs_0 ? 7'h45 : _GEN_80; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_82 = 10'h52 == io_inputs_0 ? 7'h44 : _GEN_81; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_83 = 10'h53 == io_inputs_0 ? 7'h43 : _GEN_82; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_84 = 10'h54 == io_inputs_0 ? 7'h42 : _GEN_83; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_85 = 10'h55 == io_inputs_0 ? 7'h41 : _GEN_84; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_86 = 10'h56 == io_inputs_0 ? 7'h40 : _GEN_85; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_87 = 10'h57 == io_inputs_0 ? 7'h3f : _GEN_86; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_88 = 10'h58 == io_inputs_0 ? 7'h3e : _GEN_87; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_89 = 10'h59 == io_inputs_0 ? 7'h3d : _GEN_88; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_90 = 10'h5a == io_inputs_0 ? 7'h3c : _GEN_89; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_91 = 10'h5b == io_inputs_0 ? 7'h3b : _GEN_90; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_92 = 10'h5c == io_inputs_0 ? 7'h3a : _GEN_91; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_93 = 10'h5d == io_inputs_0 ? 7'h39 : _GEN_92; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_94 = 10'h5e == io_inputs_0 ? 7'h38 : _GEN_93; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_95 = 10'h5f == io_inputs_0 ? 7'h37 : _GEN_94; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_96 = 10'h60 == io_inputs_0 ? 7'h36 : _GEN_95; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_97 = 10'h61 == io_inputs_0 ? 7'h35 : _GEN_96; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_98 = 10'h62 == io_inputs_0 ? 7'h34 : _GEN_97; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_99 = 10'h63 == io_inputs_0 ? 7'h33 : _GEN_98; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_100 = 10'h64 == io_inputs_0 ? 7'h32 : _GEN_99; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_101 = 10'h65 == io_inputs_0 ? 7'h31 : _GEN_100; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_102 = 10'h66 == io_inputs_0 ? 7'h30 : _GEN_101; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_103 = 10'h67 == io_inputs_0 ? 7'h2f : _GEN_102; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_104 = 10'h68 == io_inputs_0 ? 7'h2e : _GEN_103; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_105 = 10'h69 == io_inputs_0 ? 7'h2d : _GEN_104; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_106 = 10'h6a == io_inputs_0 ? 7'h2c : _GEN_105; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_107 = 10'h6b == io_inputs_0 ? 7'h2b : _GEN_106; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_108 = 10'h6c == io_inputs_0 ? 7'h2a : _GEN_107; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_109 = 10'h6d == io_inputs_0 ? 7'h29 : _GEN_108; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_110 = 10'h6e == io_inputs_0 ? 7'h28 : _GEN_109; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_111 = 10'h6f == io_inputs_0 ? 7'h27 : _GEN_110; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_112 = 10'h70 == io_inputs_0 ? 7'h26 : _GEN_111; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_113 = 10'h71 == io_inputs_0 ? 7'h25 : _GEN_112; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_114 = 10'h72 == io_inputs_0 ? 7'h24 : _GEN_113; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_115 = 10'h73 == io_inputs_0 ? 7'h23 : _GEN_114; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_116 = 10'h74 == io_inputs_0 ? 7'h22 : _GEN_115; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_117 = 10'h75 == io_inputs_0 ? 7'h21 : _GEN_116; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_118 = 10'h76 == io_inputs_0 ? 7'h20 : _GEN_117; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_119 = 10'h77 == io_inputs_0 ? 7'h1f : _GEN_118; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_120 = 10'h78 == io_inputs_0 ? 7'h1e : _GEN_119; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_121 = 10'h79 == io_inputs_0 ? 7'h1d : _GEN_120; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_122 = 10'h7a == io_inputs_0 ? 7'h1c : _GEN_121; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_123 = 10'h7b == io_inputs_0 ? 7'h1b : _GEN_122; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_124 = 10'h7c == io_inputs_0 ? 7'h1a : _GEN_123; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_125 = 10'h7d == io_inputs_0 ? 7'h19 : _GEN_124; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_126 = 10'h7e == io_inputs_0 ? 7'h18 : _GEN_125; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_127 = 10'h7f == io_inputs_0 ? 7'h17 : _GEN_126; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_128 = 10'h80 == io_inputs_0 ? 7'h16 : _GEN_127; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_129 = 10'h81 == io_inputs_0 ? 7'h15 : _GEN_128; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_130 = 10'h82 == io_inputs_0 ? 7'h14 : _GEN_129; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_131 = 10'h83 == io_inputs_0 ? 7'h13 : _GEN_130; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_132 = 10'h84 == io_inputs_0 ? 7'h12 : _GEN_131; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_133 = 10'h85 == io_inputs_0 ? 7'h11 : _GEN_132; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_134 = 10'h86 == io_inputs_0 ? 7'h10 : _GEN_133; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_135 = 10'h87 == io_inputs_0 ? 7'hf : _GEN_134; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_136 = 10'h88 == io_inputs_0 ? 7'he : _GEN_135; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_137 = 10'h89 == io_inputs_0 ? 7'hd : _GEN_136; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_138 = 10'h8a == io_inputs_0 ? 7'hc : _GEN_137; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_139 = 10'h8b == io_inputs_0 ? 7'hb : _GEN_138; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_140 = 10'h8c == io_inputs_0 ? 7'ha : _GEN_139; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_141 = 10'h8d == io_inputs_0 ? 7'h9 : _GEN_140; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_142 = 10'h8e == io_inputs_0 ? 7'h8 : _GEN_141; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_143 = 10'h8f == io_inputs_0 ? 7'h7 : _GEN_142; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_144 = 10'h90 == io_inputs_0 ? 7'h6 : _GEN_143; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_145 = 10'h91 == io_inputs_0 ? 7'h5 : _GEN_144; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_146 = 10'h92 == io_inputs_0 ? 7'h4 : _GEN_145; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_147 = 10'h93 == io_inputs_0 ? 7'h3 : _GEN_146; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_148 = 10'h94 == io_inputs_0 ? 7'h2 : _GEN_147; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_149 = 10'h95 == io_inputs_0 ? 7'h1 : _GEN_148; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_150 = 10'h96 == io_inputs_0 ? 7'h0 : _GEN_149; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_151 = 10'h97 == io_inputs_0 ? 7'h0 : _GEN_150; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_152 = 10'h98 == io_inputs_0 ? 7'h0 : _GEN_151; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_153 = 10'h99 == io_inputs_0 ? 7'h0 : _GEN_152; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_154 = 10'h9a == io_inputs_0 ? 7'h0 : _GEN_153; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_155 = 10'h9b == io_inputs_0 ? 7'h0 : _GEN_154; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_156 = 10'h9c == io_inputs_0 ? 7'h0 : _GEN_155; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_157 = 10'h9d == io_inputs_0 ? 7'h0 : _GEN_156; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_158 = 10'h9e == io_inputs_0 ? 7'h0 : _GEN_157; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_159 = 10'h9f == io_inputs_0 ? 7'h0 : _GEN_158; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_160 = 10'ha0 == io_inputs_0 ? 7'h0 : _GEN_159; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_161 = 10'ha1 == io_inputs_0 ? 7'h0 : _GEN_160; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_162 = 10'ha2 == io_inputs_0 ? 7'h0 : _GEN_161; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_163 = 10'ha3 == io_inputs_0 ? 7'h0 : _GEN_162; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_164 = 10'ha4 == io_inputs_0 ? 7'h0 : _GEN_163; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_165 = 10'ha5 == io_inputs_0 ? 7'h0 : _GEN_164; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_166 = 10'ha6 == io_inputs_0 ? 7'h0 : _GEN_165; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_167 = 10'ha7 == io_inputs_0 ? 7'h0 : _GEN_166; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_168 = 10'ha8 == io_inputs_0 ? 7'h0 : _GEN_167; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_169 = 10'ha9 == io_inputs_0 ? 7'h0 : _GEN_168; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_170 = 10'haa == io_inputs_0 ? 7'h0 : _GEN_169; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_171 = 10'hab == io_inputs_0 ? 7'h0 : _GEN_170; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_172 = 10'hac == io_inputs_0 ? 7'h0 : _GEN_171; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_173 = 10'had == io_inputs_0 ? 7'h0 : _GEN_172; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_174 = 10'hae == io_inputs_0 ? 7'h0 : _GEN_173; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_175 = 10'haf == io_inputs_0 ? 7'h0 : _GEN_174; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_176 = 10'hb0 == io_inputs_0 ? 7'h0 : _GEN_175; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_177 = 10'hb1 == io_inputs_0 ? 7'h0 : _GEN_176; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_178 = 10'hb2 == io_inputs_0 ? 7'h0 : _GEN_177; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_179 = 10'hb3 == io_inputs_0 ? 7'h0 : _GEN_178; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_180 = 10'hb4 == io_inputs_0 ? 7'h0 : _GEN_179; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_181 = 10'hb5 == io_inputs_0 ? 7'h0 : _GEN_180; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_182 = 10'hb6 == io_inputs_0 ? 7'h0 : _GEN_181; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_183 = 10'hb7 == io_inputs_0 ? 7'h0 : _GEN_182; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_184 = 10'hb8 == io_inputs_0 ? 7'h0 : _GEN_183; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_185 = 10'hb9 == io_inputs_0 ? 7'h0 : _GEN_184; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_186 = 10'hba == io_inputs_0 ? 7'h0 : _GEN_185; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_187 = 10'hbb == io_inputs_0 ? 7'h0 : _GEN_186; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_188 = 10'hbc == io_inputs_0 ? 7'h0 : _GEN_187; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_189 = 10'hbd == io_inputs_0 ? 7'h0 : _GEN_188; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_190 = 10'hbe == io_inputs_0 ? 7'h0 : _GEN_189; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_191 = 10'hbf == io_inputs_0 ? 7'h0 : _GEN_190; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_192 = 10'hc0 == io_inputs_0 ? 7'h0 : _GEN_191; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_193 = 10'hc1 == io_inputs_0 ? 7'h0 : _GEN_192; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_194 = 10'hc2 == io_inputs_0 ? 7'h0 : _GEN_193; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_195 = 10'hc3 == io_inputs_0 ? 7'h0 : _GEN_194; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_196 = 10'hc4 == io_inputs_0 ? 7'h0 : _GEN_195; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_197 = 10'hc5 == io_inputs_0 ? 7'h0 : _GEN_196; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_198 = 10'hc6 == io_inputs_0 ? 7'h0 : _GEN_197; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_199 = 10'hc7 == io_inputs_0 ? 7'h0 : _GEN_198; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_200 = 10'hc8 == io_inputs_0 ? 7'h0 : _GEN_199; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_201 = 10'hc9 == io_inputs_0 ? 7'h0 : _GEN_200; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_202 = 10'hca == io_inputs_0 ? 7'h0 : _GEN_201; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_203 = 10'hcb == io_inputs_0 ? 7'h0 : _GEN_202; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_204 = 10'hcc == io_inputs_0 ? 7'h0 : _GEN_203; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_205 = 10'hcd == io_inputs_0 ? 7'h0 : _GEN_204; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_206 = 10'hce == io_inputs_0 ? 7'h0 : _GEN_205; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_207 = 10'hcf == io_inputs_0 ? 7'h0 : _GEN_206; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_208 = 10'hd0 == io_inputs_0 ? 7'h0 : _GEN_207; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_209 = 10'hd1 == io_inputs_0 ? 7'h0 : _GEN_208; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_210 = 10'hd2 == io_inputs_0 ? 7'h0 : _GEN_209; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_211 = 10'hd3 == io_inputs_0 ? 7'h0 : _GEN_210; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_212 = 10'hd4 == io_inputs_0 ? 7'h0 : _GEN_211; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_213 = 10'hd5 == io_inputs_0 ? 7'h0 : _GEN_212; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_214 = 10'hd6 == io_inputs_0 ? 7'h0 : _GEN_213; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_215 = 10'hd7 == io_inputs_0 ? 7'h0 : _GEN_214; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_216 = 10'hd8 == io_inputs_0 ? 7'h0 : _GEN_215; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_217 = 10'hd9 == io_inputs_0 ? 7'h0 : _GEN_216; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_218 = 10'hda == io_inputs_0 ? 7'h0 : _GEN_217; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_219 = 10'hdb == io_inputs_0 ? 7'h0 : _GEN_218; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_220 = 10'hdc == io_inputs_0 ? 7'h0 : _GEN_219; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_221 = 10'hdd == io_inputs_0 ? 7'h0 : _GEN_220; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_222 = 10'hde == io_inputs_0 ? 7'h0 : _GEN_221; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_223 = 10'hdf == io_inputs_0 ? 7'h0 : _GEN_222; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_224 = 10'he0 == io_inputs_0 ? 7'h0 : _GEN_223; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_225 = 10'he1 == io_inputs_0 ? 7'h0 : _GEN_224; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_226 = 10'he2 == io_inputs_0 ? 7'h0 : _GEN_225; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_227 = 10'he3 == io_inputs_0 ? 7'h0 : _GEN_226; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_228 = 10'he4 == io_inputs_0 ? 7'h0 : _GEN_227; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_229 = 10'he5 == io_inputs_0 ? 7'h0 : _GEN_228; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_230 = 10'he6 == io_inputs_0 ? 7'h0 : _GEN_229; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_231 = 10'he7 == io_inputs_0 ? 7'h0 : _GEN_230; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_232 = 10'he8 == io_inputs_0 ? 7'h0 : _GEN_231; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_233 = 10'he9 == io_inputs_0 ? 7'h0 : _GEN_232; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_234 = 10'hea == io_inputs_0 ? 7'h0 : _GEN_233; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_235 = 10'heb == io_inputs_0 ? 7'h0 : _GEN_234; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_236 = 10'hec == io_inputs_0 ? 7'h0 : _GEN_235; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_237 = 10'hed == io_inputs_0 ? 7'h0 : _GEN_236; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_238 = 10'hee == io_inputs_0 ? 7'h0 : _GEN_237; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_239 = 10'hef == io_inputs_0 ? 7'h0 : _GEN_238; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_240 = 10'hf0 == io_inputs_0 ? 7'h0 : _GEN_239; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_241 = 10'hf1 == io_inputs_0 ? 7'h0 : _GEN_240; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_242 = 10'hf2 == io_inputs_0 ? 7'h0 : _GEN_241; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_243 = 10'hf3 == io_inputs_0 ? 7'h0 : _GEN_242; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_244 = 10'hf4 == io_inputs_0 ? 7'h0 : _GEN_243; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_245 = 10'hf5 == io_inputs_0 ? 7'h0 : _GEN_244; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_246 = 10'hf6 == io_inputs_0 ? 7'h0 : _GEN_245; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_247 = 10'hf7 == io_inputs_0 ? 7'h0 : _GEN_246; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_248 = 10'hf8 == io_inputs_0 ? 7'h0 : _GEN_247; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_249 = 10'hf9 == io_inputs_0 ? 7'h0 : _GEN_248; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_250 = 10'hfa == io_inputs_0 ? 7'h0 : _GEN_249; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_251 = 10'hfb == io_inputs_0 ? 7'h0 : _GEN_250; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_252 = 10'hfc == io_inputs_0 ? 7'h0 : _GEN_251; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_253 = 10'hfd == io_inputs_0 ? 7'h0 : _GEN_252; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_254 = 10'hfe == io_inputs_0 ? 7'h0 : _GEN_253; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_255 = 10'hff == io_inputs_0 ? 7'h0 : _GEN_254; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_256 = 10'h100 == io_inputs_0 ? 7'h0 : _GEN_255; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_257 = 10'h101 == io_inputs_0 ? 7'h0 : _GEN_256; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_258 = 10'h102 == io_inputs_0 ? 7'h0 : _GEN_257; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_259 = 10'h103 == io_inputs_0 ? 7'h0 : _GEN_258; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_260 = 10'h104 == io_inputs_0 ? 7'h0 : _GEN_259; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_261 = 10'h105 == io_inputs_0 ? 7'h0 : _GEN_260; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_262 = 10'h106 == io_inputs_0 ? 7'h0 : _GEN_261; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_263 = 10'h107 == io_inputs_0 ? 7'h0 : _GEN_262; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_264 = 10'h108 == io_inputs_0 ? 7'h0 : _GEN_263; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_265 = 10'h109 == io_inputs_0 ? 7'h0 : _GEN_264; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_266 = 10'h10a == io_inputs_0 ? 7'h0 : _GEN_265; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_267 = 10'h10b == io_inputs_0 ? 7'h0 : _GEN_266; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_268 = 10'h10c == io_inputs_0 ? 7'h0 : _GEN_267; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_269 = 10'h10d == io_inputs_0 ? 7'h0 : _GEN_268; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_270 = 10'h10e == io_inputs_0 ? 7'h0 : _GEN_269; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_271 = 10'h10f == io_inputs_0 ? 7'h0 : _GEN_270; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_272 = 10'h110 == io_inputs_0 ? 7'h0 : _GEN_271; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_273 = 10'h111 == io_inputs_0 ? 7'h0 : _GEN_272; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_274 = 10'h112 == io_inputs_0 ? 7'h0 : _GEN_273; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_275 = 10'h113 == io_inputs_0 ? 7'h0 : _GEN_274; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_276 = 10'h114 == io_inputs_0 ? 7'h0 : _GEN_275; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_277 = 10'h115 == io_inputs_0 ? 7'h0 : _GEN_276; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_278 = 10'h116 == io_inputs_0 ? 7'h0 : _GEN_277; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_279 = 10'h117 == io_inputs_0 ? 7'h0 : _GEN_278; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_280 = 10'h118 == io_inputs_0 ? 7'h0 : _GEN_279; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_281 = 10'h119 == io_inputs_0 ? 7'h0 : _GEN_280; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_282 = 10'h11a == io_inputs_0 ? 7'h0 : _GEN_281; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_283 = 10'h11b == io_inputs_0 ? 7'h0 : _GEN_282; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_284 = 10'h11c == io_inputs_0 ? 7'h0 : _GEN_283; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_285 = 10'h11d == io_inputs_0 ? 7'h0 : _GEN_284; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_286 = 10'h11e == io_inputs_0 ? 7'h0 : _GEN_285; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_287 = 10'h11f == io_inputs_0 ? 7'h0 : _GEN_286; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_288 = 10'h120 == io_inputs_0 ? 7'h0 : _GEN_287; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_289 = 10'h121 == io_inputs_0 ? 7'h0 : _GEN_288; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_290 = 10'h122 == io_inputs_0 ? 7'h0 : _GEN_289; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_291 = 10'h123 == io_inputs_0 ? 7'h0 : _GEN_290; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_292 = 10'h124 == io_inputs_0 ? 7'h0 : _GEN_291; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_293 = 10'h125 == io_inputs_0 ? 7'h0 : _GEN_292; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_294 = 10'h126 == io_inputs_0 ? 7'h0 : _GEN_293; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_295 = 10'h127 == io_inputs_0 ? 7'h0 : _GEN_294; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_296 = 10'h128 == io_inputs_0 ? 7'h0 : _GEN_295; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_297 = 10'h129 == io_inputs_0 ? 7'h0 : _GEN_296; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_298 = 10'h12a == io_inputs_0 ? 7'h0 : _GEN_297; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_299 = 10'h12b == io_inputs_0 ? 7'h0 : _GEN_298; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_300 = 10'h12c == io_inputs_0 ? 7'h0 : _GEN_299; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_301 = 10'h12d == io_inputs_0 ? 7'h0 : _GEN_300; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_302 = 10'h12e == io_inputs_0 ? 7'h0 : _GEN_301; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_303 = 10'h12f == io_inputs_0 ? 7'h0 : _GEN_302; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_304 = 10'h130 == io_inputs_0 ? 7'h0 : _GEN_303; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_305 = 10'h131 == io_inputs_0 ? 7'h0 : _GEN_304; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_306 = 10'h132 == io_inputs_0 ? 7'h0 : _GEN_305; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_307 = 10'h133 == io_inputs_0 ? 7'h0 : _GEN_306; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_308 = 10'h134 == io_inputs_0 ? 7'h0 : _GEN_307; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_309 = 10'h135 == io_inputs_0 ? 7'h0 : _GEN_308; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_310 = 10'h136 == io_inputs_0 ? 7'h0 : _GEN_309; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_311 = 10'h137 == io_inputs_0 ? 7'h0 : _GEN_310; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_312 = 10'h138 == io_inputs_0 ? 7'h0 : _GEN_311; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_313 = 10'h139 == io_inputs_0 ? 7'h0 : _GEN_312; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_314 = 10'h13a == io_inputs_0 ? 7'h0 : _GEN_313; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_315 = 10'h13b == io_inputs_0 ? 7'h0 : _GEN_314; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_316 = 10'h13c == io_inputs_0 ? 7'h0 : _GEN_315; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_317 = 10'h13d == io_inputs_0 ? 7'h0 : _GEN_316; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_318 = 10'h13e == io_inputs_0 ? 7'h0 : _GEN_317; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_319 = 10'h13f == io_inputs_0 ? 7'h0 : _GEN_318; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_320 = 10'h140 == io_inputs_0 ? 7'h0 : _GEN_319; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_321 = 10'h141 == io_inputs_0 ? 7'h0 : _GEN_320; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_322 = 10'h142 == io_inputs_0 ? 7'h0 : _GEN_321; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_323 = 10'h143 == io_inputs_0 ? 7'h0 : _GEN_322; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_324 = 10'h144 == io_inputs_0 ? 7'h0 : _GEN_323; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_325 = 10'h145 == io_inputs_0 ? 7'h0 : _GEN_324; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_326 = 10'h146 == io_inputs_0 ? 7'h0 : _GEN_325; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_327 = 10'h147 == io_inputs_0 ? 7'h0 : _GEN_326; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_328 = 10'h148 == io_inputs_0 ? 7'h0 : _GEN_327; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_329 = 10'h149 == io_inputs_0 ? 7'h0 : _GEN_328; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_330 = 10'h14a == io_inputs_0 ? 7'h0 : _GEN_329; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_331 = 10'h14b == io_inputs_0 ? 7'h0 : _GEN_330; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_332 = 10'h14c == io_inputs_0 ? 7'h0 : _GEN_331; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_333 = 10'h14d == io_inputs_0 ? 7'h0 : _GEN_332; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_334 = 10'h14e == io_inputs_0 ? 7'h0 : _GEN_333; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_335 = 10'h14f == io_inputs_0 ? 7'h0 : _GEN_334; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_336 = 10'h150 == io_inputs_0 ? 7'h0 : _GEN_335; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_337 = 10'h151 == io_inputs_0 ? 7'h0 : _GEN_336; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_338 = 10'h152 == io_inputs_0 ? 7'h0 : _GEN_337; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_339 = 10'h153 == io_inputs_0 ? 7'h0 : _GEN_338; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_340 = 10'h154 == io_inputs_0 ? 7'h0 : _GEN_339; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_341 = 10'h155 == io_inputs_0 ? 7'h0 : _GEN_340; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_342 = 10'h156 == io_inputs_0 ? 7'h0 : _GEN_341; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_343 = 10'h157 == io_inputs_0 ? 7'h0 : _GEN_342; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_344 = 10'h158 == io_inputs_0 ? 7'h0 : _GEN_343; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_345 = 10'h159 == io_inputs_0 ? 7'h0 : _GEN_344; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_346 = 10'h15a == io_inputs_0 ? 7'h0 : _GEN_345; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_347 = 10'h15b == io_inputs_0 ? 7'h0 : _GEN_346; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_348 = 10'h15c == io_inputs_0 ? 7'h0 : _GEN_347; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_349 = 10'h15d == io_inputs_0 ? 7'h0 : _GEN_348; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_350 = 10'h15e == io_inputs_0 ? 7'h0 : _GEN_349; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_351 = 10'h15f == io_inputs_0 ? 7'h0 : _GEN_350; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_352 = 10'h160 == io_inputs_0 ? 7'h0 : _GEN_351; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_353 = 10'h161 == io_inputs_0 ? 7'h0 : _GEN_352; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_354 = 10'h162 == io_inputs_0 ? 7'h0 : _GEN_353; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_355 = 10'h163 == io_inputs_0 ? 7'h0 : _GEN_354; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_356 = 10'h164 == io_inputs_0 ? 7'h0 : _GEN_355; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_357 = 10'h165 == io_inputs_0 ? 7'h0 : _GEN_356; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_358 = 10'h166 == io_inputs_0 ? 7'h0 : _GEN_357; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_359 = 10'h167 == io_inputs_0 ? 7'h0 : _GEN_358; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_360 = 10'h168 == io_inputs_0 ? 7'h0 : _GEN_359; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_361 = 10'h169 == io_inputs_0 ? 7'h0 : _GEN_360; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_362 = 10'h16a == io_inputs_0 ? 7'h0 : _GEN_361; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_363 = 10'h16b == io_inputs_0 ? 7'h0 : _GEN_362; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_364 = 10'h16c == io_inputs_0 ? 7'h0 : _GEN_363; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_365 = 10'h16d == io_inputs_0 ? 7'h0 : _GEN_364; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_366 = 10'h16e == io_inputs_0 ? 7'h0 : _GEN_365; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_367 = 10'h16f == io_inputs_0 ? 7'h0 : _GEN_366; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_368 = 10'h170 == io_inputs_0 ? 7'h0 : _GEN_367; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_369 = 10'h171 == io_inputs_0 ? 7'h0 : _GEN_368; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_370 = 10'h172 == io_inputs_0 ? 7'h0 : _GEN_369; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_371 = 10'h173 == io_inputs_0 ? 7'h0 : _GEN_370; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_372 = 10'h174 == io_inputs_0 ? 7'h0 : _GEN_371; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_373 = 10'h175 == io_inputs_0 ? 7'h0 : _GEN_372; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_374 = 10'h176 == io_inputs_0 ? 7'h0 : _GEN_373; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_375 = 10'h177 == io_inputs_0 ? 7'h0 : _GEN_374; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_376 = 10'h178 == io_inputs_0 ? 7'h0 : _GEN_375; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_377 = 10'h179 == io_inputs_0 ? 7'h0 : _GEN_376; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_378 = 10'h17a == io_inputs_0 ? 7'h0 : _GEN_377; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_379 = 10'h17b == io_inputs_0 ? 7'h0 : _GEN_378; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_380 = 10'h17c == io_inputs_0 ? 7'h0 : _GEN_379; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_381 = 10'h17d == io_inputs_0 ? 7'h0 : _GEN_380; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_382 = 10'h17e == io_inputs_0 ? 7'h0 : _GEN_381; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_383 = 10'h17f == io_inputs_0 ? 7'h0 : _GEN_382; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_384 = 10'h180 == io_inputs_0 ? 7'h0 : _GEN_383; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_385 = 10'h181 == io_inputs_0 ? 7'h0 : _GEN_384; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_386 = 10'h182 == io_inputs_0 ? 7'h0 : _GEN_385; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_387 = 10'h183 == io_inputs_0 ? 7'h0 : _GEN_386; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_388 = 10'h184 == io_inputs_0 ? 7'h0 : _GEN_387; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_389 = 10'h185 == io_inputs_0 ? 7'h0 : _GEN_388; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_390 = 10'h186 == io_inputs_0 ? 7'h0 : _GEN_389; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_391 = 10'h187 == io_inputs_0 ? 7'h0 : _GEN_390; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_392 = 10'h188 == io_inputs_0 ? 7'h0 : _GEN_391; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_393 = 10'h189 == io_inputs_0 ? 7'h0 : _GEN_392; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_394 = 10'h18a == io_inputs_0 ? 7'h0 : _GEN_393; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_395 = 10'h18b == io_inputs_0 ? 7'h0 : _GEN_394; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_396 = 10'h18c == io_inputs_0 ? 7'h0 : _GEN_395; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_397 = 10'h18d == io_inputs_0 ? 7'h0 : _GEN_396; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_398 = 10'h18e == io_inputs_0 ? 7'h0 : _GEN_397; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_399 = 10'h18f == io_inputs_0 ? 7'h0 : _GEN_398; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_400 = 10'h190 == io_inputs_0 ? 7'h0 : _GEN_399; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_401 = 10'h191 == io_inputs_0 ? 7'h0 : _GEN_400; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_402 = 10'h192 == io_inputs_0 ? 7'h0 : _GEN_401; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_403 = 10'h193 == io_inputs_0 ? 7'h0 : _GEN_402; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_404 = 10'h194 == io_inputs_0 ? 7'h0 : _GEN_403; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_405 = 10'h195 == io_inputs_0 ? 7'h0 : _GEN_404; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_406 = 10'h196 == io_inputs_0 ? 7'h0 : _GEN_405; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_407 = 10'h197 == io_inputs_0 ? 7'h0 : _GEN_406; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_408 = 10'h198 == io_inputs_0 ? 7'h0 : _GEN_407; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_409 = 10'h199 == io_inputs_0 ? 7'h0 : _GEN_408; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_410 = 10'h19a == io_inputs_0 ? 7'h0 : _GEN_409; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_411 = 10'h19b == io_inputs_0 ? 7'h0 : _GEN_410; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_412 = 10'h19c == io_inputs_0 ? 7'h0 : _GEN_411; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_413 = 10'h19d == io_inputs_0 ? 7'h0 : _GEN_412; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_414 = 10'h19e == io_inputs_0 ? 7'h0 : _GEN_413; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_415 = 10'h19f == io_inputs_0 ? 7'h0 : _GEN_414; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_416 = 10'h1a0 == io_inputs_0 ? 7'h0 : _GEN_415; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_417 = 10'h1a1 == io_inputs_0 ? 7'h0 : _GEN_416; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_418 = 10'h1a2 == io_inputs_0 ? 7'h0 : _GEN_417; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_419 = 10'h1a3 == io_inputs_0 ? 7'h0 : _GEN_418; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_420 = 10'h1a4 == io_inputs_0 ? 7'h0 : _GEN_419; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_421 = 10'h1a5 == io_inputs_0 ? 7'h0 : _GEN_420; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_422 = 10'h1a6 == io_inputs_0 ? 7'h0 : _GEN_421; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_423 = 10'h1a7 == io_inputs_0 ? 7'h0 : _GEN_422; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_424 = 10'h1a8 == io_inputs_0 ? 7'h0 : _GEN_423; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_425 = 10'h1a9 == io_inputs_0 ? 7'h0 : _GEN_424; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_426 = 10'h1aa == io_inputs_0 ? 7'h0 : _GEN_425; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_427 = 10'h1ab == io_inputs_0 ? 7'h0 : _GEN_426; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_428 = 10'h1ac == io_inputs_0 ? 7'h0 : _GEN_427; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_429 = 10'h1ad == io_inputs_0 ? 7'h0 : _GEN_428; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_430 = 10'h1ae == io_inputs_0 ? 7'h0 : _GEN_429; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_431 = 10'h1af == io_inputs_0 ? 7'h0 : _GEN_430; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_432 = 10'h1b0 == io_inputs_0 ? 7'h0 : _GEN_431; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_433 = 10'h1b1 == io_inputs_0 ? 7'h0 : _GEN_432; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_434 = 10'h1b2 == io_inputs_0 ? 7'h0 : _GEN_433; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_435 = 10'h1b3 == io_inputs_0 ? 7'h0 : _GEN_434; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_436 = 10'h1b4 == io_inputs_0 ? 7'h0 : _GEN_435; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_437 = 10'h1b5 == io_inputs_0 ? 7'h0 : _GEN_436; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_438 = 10'h1b6 == io_inputs_0 ? 7'h0 : _GEN_437; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_439 = 10'h1b7 == io_inputs_0 ? 7'h0 : _GEN_438; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_440 = 10'h1b8 == io_inputs_0 ? 7'h0 : _GEN_439; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_441 = 10'h1b9 == io_inputs_0 ? 7'h0 : _GEN_440; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_442 = 10'h1ba == io_inputs_0 ? 7'h0 : _GEN_441; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_443 = 10'h1bb == io_inputs_0 ? 7'h0 : _GEN_442; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_444 = 10'h1bc == io_inputs_0 ? 7'h0 : _GEN_443; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_445 = 10'h1bd == io_inputs_0 ? 7'h0 : _GEN_444; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_446 = 10'h1be == io_inputs_0 ? 7'h0 : _GEN_445; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_447 = 10'h1bf == io_inputs_0 ? 7'h0 : _GEN_446; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_448 = 10'h1c0 == io_inputs_0 ? 7'h0 : _GEN_447; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_449 = 10'h1c1 == io_inputs_0 ? 7'h0 : _GEN_448; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_450 = 10'h1c2 == io_inputs_0 ? 7'h0 : _GEN_449; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_451 = 10'h1c3 == io_inputs_0 ? 7'h0 : _GEN_450; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_452 = 10'h1c4 == io_inputs_0 ? 7'h0 : _GEN_451; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_453 = 10'h1c5 == io_inputs_0 ? 7'h0 : _GEN_452; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_454 = 10'h1c6 == io_inputs_0 ? 7'h0 : _GEN_453; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_455 = 10'h1c7 == io_inputs_0 ? 7'h0 : _GEN_454; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_456 = 10'h1c8 == io_inputs_0 ? 7'h0 : _GEN_455; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_457 = 10'h1c9 == io_inputs_0 ? 7'h0 : _GEN_456; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_458 = 10'h1ca == io_inputs_0 ? 7'h0 : _GEN_457; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_459 = 10'h1cb == io_inputs_0 ? 7'h0 : _GEN_458; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_460 = 10'h1cc == io_inputs_0 ? 7'h0 : _GEN_459; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_461 = 10'h1cd == io_inputs_0 ? 7'h0 : _GEN_460; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_462 = 10'h1ce == io_inputs_0 ? 7'h0 : _GEN_461; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_463 = 10'h1cf == io_inputs_0 ? 7'h0 : _GEN_462; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_464 = 10'h1d0 == io_inputs_0 ? 7'h0 : _GEN_463; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_465 = 10'h1d1 == io_inputs_0 ? 7'h0 : _GEN_464; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_466 = 10'h1d2 == io_inputs_0 ? 7'h0 : _GEN_465; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_467 = 10'h1d3 == io_inputs_0 ? 7'h0 : _GEN_466; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_468 = 10'h1d4 == io_inputs_0 ? 7'h0 : _GEN_467; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_469 = 10'h1d5 == io_inputs_0 ? 7'h0 : _GEN_468; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_470 = 10'h1d6 == io_inputs_0 ? 7'h0 : _GEN_469; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_471 = 10'h1d7 == io_inputs_0 ? 7'h0 : _GEN_470; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_472 = 10'h1d8 == io_inputs_0 ? 7'h0 : _GEN_471; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_473 = 10'h1d9 == io_inputs_0 ? 7'h0 : _GEN_472; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_474 = 10'h1da == io_inputs_0 ? 7'h0 : _GEN_473; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_475 = 10'h1db == io_inputs_0 ? 7'h0 : _GEN_474; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_476 = 10'h1dc == io_inputs_0 ? 7'h0 : _GEN_475; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_477 = 10'h1dd == io_inputs_0 ? 7'h0 : _GEN_476; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_478 = 10'h1de == io_inputs_0 ? 7'h0 : _GEN_477; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_479 = 10'h1df == io_inputs_0 ? 7'h0 : _GEN_478; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_480 = 10'h1e0 == io_inputs_0 ? 7'h0 : _GEN_479; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_481 = 10'h1e1 == io_inputs_0 ? 7'h0 : _GEN_480; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_482 = 10'h1e2 == io_inputs_0 ? 7'h0 : _GEN_481; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_483 = 10'h1e3 == io_inputs_0 ? 7'h0 : _GEN_482; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_484 = 10'h1e4 == io_inputs_0 ? 7'h0 : _GEN_483; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_485 = 10'h1e5 == io_inputs_0 ? 7'h0 : _GEN_484; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_486 = 10'h1e6 == io_inputs_0 ? 7'h0 : _GEN_485; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_487 = 10'h1e7 == io_inputs_0 ? 7'h0 : _GEN_486; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_488 = 10'h1e8 == io_inputs_0 ? 7'h0 : _GEN_487; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_489 = 10'h1e9 == io_inputs_0 ? 7'h0 : _GEN_488; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_490 = 10'h1ea == io_inputs_0 ? 7'h0 : _GEN_489; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_491 = 10'h1eb == io_inputs_0 ? 7'h0 : _GEN_490; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_492 = 10'h1ec == io_inputs_0 ? 7'h0 : _GEN_491; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_493 = 10'h1ed == io_inputs_0 ? 7'h0 : _GEN_492; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_494 = 10'h1ee == io_inputs_0 ? 7'h0 : _GEN_493; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_495 = 10'h1ef == io_inputs_0 ? 7'h0 : _GEN_494; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_496 = 10'h1f0 == io_inputs_0 ? 7'h0 : _GEN_495; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_497 = 10'h1f1 == io_inputs_0 ? 7'h0 : _GEN_496; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_498 = 10'h1f2 == io_inputs_0 ? 7'h0 : _GEN_497; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_499 = 10'h1f3 == io_inputs_0 ? 7'h0 : _GEN_498; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_500 = 10'h1f4 == io_inputs_0 ? 7'h0 : _GEN_499; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_501 = 10'h1f5 == io_inputs_0 ? 7'h0 : _GEN_500; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_502 = 10'h1f6 == io_inputs_0 ? 7'h0 : _GEN_501; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_503 = 10'h1f7 == io_inputs_0 ? 7'h0 : _GEN_502; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_504 = 10'h1f8 == io_inputs_0 ? 7'h0 : _GEN_503; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_505 = 10'h1f9 == io_inputs_0 ? 7'h0 : _GEN_504; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_506 = 10'h1fa == io_inputs_0 ? 7'h0 : _GEN_505; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_507 = 10'h1fb == io_inputs_0 ? 7'h0 : _GEN_506; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_508 = 10'h1fc == io_inputs_0 ? 7'h0 : _GEN_507; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_509 = 10'h1fd == io_inputs_0 ? 7'h0 : _GEN_508; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_510 = 10'h1fe == io_inputs_0 ? 7'h0 : _GEN_509; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_511 = 10'h1ff == io_inputs_0 ? 7'h0 : _GEN_510; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_512 = 10'h200 == io_inputs_0 ? 7'h0 : _GEN_511; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_513 = 10'h201 == io_inputs_0 ? 7'h0 : _GEN_512; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_514 = 10'h202 == io_inputs_0 ? 7'h0 : _GEN_513; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_515 = 10'h203 == io_inputs_0 ? 7'h0 : _GEN_514; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_516 = 10'h204 == io_inputs_0 ? 7'h0 : _GEN_515; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_517 = 10'h205 == io_inputs_0 ? 7'h0 : _GEN_516; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_518 = 10'h206 == io_inputs_0 ? 7'h0 : _GEN_517; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_519 = 10'h207 == io_inputs_0 ? 7'h0 : _GEN_518; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_520 = 10'h208 == io_inputs_0 ? 7'h0 : _GEN_519; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_521 = 10'h209 == io_inputs_0 ? 7'h0 : _GEN_520; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_522 = 10'h20a == io_inputs_0 ? 7'h0 : _GEN_521; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_523 = 10'h20b == io_inputs_0 ? 7'h0 : _GEN_522; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_524 = 10'h20c == io_inputs_0 ? 7'h0 : _GEN_523; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_525 = 10'h20d == io_inputs_0 ? 7'h0 : _GEN_524; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_526 = 10'h20e == io_inputs_0 ? 7'h0 : _GEN_525; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_527 = 10'h20f == io_inputs_0 ? 7'h0 : _GEN_526; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_528 = 10'h210 == io_inputs_0 ? 7'h0 : _GEN_527; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_529 = 10'h211 == io_inputs_0 ? 7'h0 : _GEN_528; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_530 = 10'h212 == io_inputs_0 ? 7'h0 : _GEN_529; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_531 = 10'h213 == io_inputs_0 ? 7'h0 : _GEN_530; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_532 = 10'h214 == io_inputs_0 ? 7'h0 : _GEN_531; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_533 = 10'h215 == io_inputs_0 ? 7'h0 : _GEN_532; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_534 = 10'h216 == io_inputs_0 ? 7'h0 : _GEN_533; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_535 = 10'h217 == io_inputs_0 ? 7'h0 : _GEN_534; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_536 = 10'h218 == io_inputs_0 ? 7'h0 : _GEN_535; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_537 = 10'h219 == io_inputs_0 ? 7'h0 : _GEN_536; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_538 = 10'h21a == io_inputs_0 ? 7'h0 : _GEN_537; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_539 = 10'h21b == io_inputs_0 ? 7'h0 : _GEN_538; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_540 = 10'h21c == io_inputs_0 ? 7'h0 : _GEN_539; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_541 = 10'h21d == io_inputs_0 ? 7'h0 : _GEN_540; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_542 = 10'h21e == io_inputs_0 ? 7'h0 : _GEN_541; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_543 = 10'h21f == io_inputs_0 ? 7'h0 : _GEN_542; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_544 = 10'h220 == io_inputs_0 ? 7'h0 : _GEN_543; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_545 = 10'h221 == io_inputs_0 ? 7'h0 : _GEN_544; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_546 = 10'h222 == io_inputs_0 ? 7'h0 : _GEN_545; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_547 = 10'h223 == io_inputs_0 ? 7'h0 : _GEN_546; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_548 = 10'h224 == io_inputs_0 ? 7'h0 : _GEN_547; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_549 = 10'h225 == io_inputs_0 ? 7'h0 : _GEN_548; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_550 = 10'h226 == io_inputs_0 ? 7'h0 : _GEN_549; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_551 = 10'h227 == io_inputs_0 ? 7'h0 : _GEN_550; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_552 = 10'h228 == io_inputs_0 ? 7'h0 : _GEN_551; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_553 = 10'h229 == io_inputs_0 ? 7'h0 : _GEN_552; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_554 = 10'h22a == io_inputs_0 ? 7'h0 : _GEN_553; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_555 = 10'h22b == io_inputs_0 ? 7'h0 : _GEN_554; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_556 = 10'h22c == io_inputs_0 ? 7'h0 : _GEN_555; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_557 = 10'h22d == io_inputs_0 ? 7'h0 : _GEN_556; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_558 = 10'h22e == io_inputs_0 ? 7'h0 : _GEN_557; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_559 = 10'h22f == io_inputs_0 ? 7'h0 : _GEN_558; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_560 = 10'h230 == io_inputs_0 ? 7'h0 : _GEN_559; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_561 = 10'h231 == io_inputs_0 ? 7'h0 : _GEN_560; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_562 = 10'h232 == io_inputs_0 ? 7'h0 : _GEN_561; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_563 = 10'h233 == io_inputs_0 ? 7'h0 : _GEN_562; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_564 = 10'h234 == io_inputs_0 ? 7'h0 : _GEN_563; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_565 = 10'h235 == io_inputs_0 ? 7'h0 : _GEN_564; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_566 = 10'h236 == io_inputs_0 ? 7'h0 : _GEN_565; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_567 = 10'h237 == io_inputs_0 ? 7'h0 : _GEN_566; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_568 = 10'h238 == io_inputs_0 ? 7'h0 : _GEN_567; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_569 = 10'h239 == io_inputs_0 ? 7'h0 : _GEN_568; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_570 = 10'h23a == io_inputs_0 ? 7'h0 : _GEN_569; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_571 = 10'h23b == io_inputs_0 ? 7'h0 : _GEN_570; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_572 = 10'h23c == io_inputs_0 ? 7'h0 : _GEN_571; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_573 = 10'h23d == io_inputs_0 ? 7'h0 : _GEN_572; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_574 = 10'h23e == io_inputs_0 ? 7'h0 : _GEN_573; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_575 = 10'h23f == io_inputs_0 ? 7'h0 : _GEN_574; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_576 = 10'h240 == io_inputs_0 ? 7'h0 : _GEN_575; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_577 = 10'h241 == io_inputs_0 ? 7'h0 : _GEN_576; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_578 = 10'h242 == io_inputs_0 ? 7'h0 : _GEN_577; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_579 = 10'h243 == io_inputs_0 ? 7'h0 : _GEN_578; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_580 = 10'h244 == io_inputs_0 ? 7'h0 : _GEN_579; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_581 = 10'h245 == io_inputs_0 ? 7'h0 : _GEN_580; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_582 = 10'h246 == io_inputs_0 ? 7'h0 : _GEN_581; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_583 = 10'h247 == io_inputs_0 ? 7'h0 : _GEN_582; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_584 = 10'h248 == io_inputs_0 ? 7'h0 : _GEN_583; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_585 = 10'h249 == io_inputs_0 ? 7'h0 : _GEN_584; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_586 = 10'h24a == io_inputs_0 ? 7'h0 : _GEN_585; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_587 = 10'h24b == io_inputs_0 ? 7'h0 : _GEN_586; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_588 = 10'h24c == io_inputs_0 ? 7'h0 : _GEN_587; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_589 = 10'h24d == io_inputs_0 ? 7'h0 : _GEN_588; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_590 = 10'h24e == io_inputs_0 ? 7'h0 : _GEN_589; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_591 = 10'h24f == io_inputs_0 ? 7'h0 : _GEN_590; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_592 = 10'h250 == io_inputs_0 ? 7'h0 : _GEN_591; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_593 = 10'h251 == io_inputs_0 ? 7'h0 : _GEN_592; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_594 = 10'h252 == io_inputs_0 ? 7'h0 : _GEN_593; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_595 = 10'h253 == io_inputs_0 ? 7'h0 : _GEN_594; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_596 = 10'h254 == io_inputs_0 ? 7'h0 : _GEN_595; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_597 = 10'h255 == io_inputs_0 ? 7'h0 : _GEN_596; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_598 = 10'h256 == io_inputs_0 ? 7'h0 : _GEN_597; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_599 = 10'h257 == io_inputs_0 ? 7'h0 : _GEN_598; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_600 = 10'h258 == io_inputs_0 ? 7'h0 : _GEN_599; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_601 = 10'h259 == io_inputs_0 ? 7'h0 : _GEN_600; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_602 = 10'h25a == io_inputs_0 ? 7'h0 : _GEN_601; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_603 = 10'h25b == io_inputs_0 ? 7'h0 : _GEN_602; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_604 = 10'h25c == io_inputs_0 ? 7'h0 : _GEN_603; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_605 = 10'h25d == io_inputs_0 ? 7'h0 : _GEN_604; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_606 = 10'h25e == io_inputs_0 ? 7'h0 : _GEN_605; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_607 = 10'h25f == io_inputs_0 ? 7'h0 : _GEN_606; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_608 = 10'h260 == io_inputs_0 ? 7'h0 : _GEN_607; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_609 = 10'h261 == io_inputs_0 ? 7'h0 : _GEN_608; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_610 = 10'h262 == io_inputs_0 ? 7'h0 : _GEN_609; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_611 = 10'h263 == io_inputs_0 ? 7'h0 : _GEN_610; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_612 = 10'h264 == io_inputs_0 ? 7'h0 : _GEN_611; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_613 = 10'h265 == io_inputs_0 ? 7'h0 : _GEN_612; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_614 = 10'h266 == io_inputs_0 ? 7'h0 : _GEN_613; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_615 = 10'h267 == io_inputs_0 ? 7'h0 : _GEN_614; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_616 = 10'h268 == io_inputs_0 ? 7'h0 : _GEN_615; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_617 = 10'h269 == io_inputs_0 ? 7'h0 : _GEN_616; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_618 = 10'h26a == io_inputs_0 ? 7'h0 : _GEN_617; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_619 = 10'h26b == io_inputs_0 ? 7'h0 : _GEN_618; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_620 = 10'h26c == io_inputs_0 ? 7'h0 : _GEN_619; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_621 = 10'h26d == io_inputs_0 ? 7'h0 : _GEN_620; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_622 = 10'h26e == io_inputs_0 ? 7'h0 : _GEN_621; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_623 = 10'h26f == io_inputs_0 ? 7'h0 : _GEN_622; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_624 = 10'h270 == io_inputs_0 ? 7'h0 : _GEN_623; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_625 = 10'h271 == io_inputs_0 ? 7'h0 : _GEN_624; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_626 = 10'h272 == io_inputs_0 ? 7'h0 : _GEN_625; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_627 = 10'h273 == io_inputs_0 ? 7'h0 : _GEN_626; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_628 = 10'h274 == io_inputs_0 ? 7'h0 : _GEN_627; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_629 = 10'h275 == io_inputs_0 ? 7'h0 : _GEN_628; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_630 = 10'h276 == io_inputs_0 ? 7'h0 : _GEN_629; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_631 = 10'h277 == io_inputs_0 ? 7'h0 : _GEN_630; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_632 = 10'h278 == io_inputs_0 ? 7'h0 : _GEN_631; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_633 = 10'h279 == io_inputs_0 ? 7'h0 : _GEN_632; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_634 = 10'h27a == io_inputs_0 ? 7'h0 : _GEN_633; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_635 = 10'h27b == io_inputs_0 ? 7'h0 : _GEN_634; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_636 = 10'h27c == io_inputs_0 ? 7'h0 : _GEN_635; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_637 = 10'h27d == io_inputs_0 ? 7'h0 : _GEN_636; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_638 = 10'h27e == io_inputs_0 ? 7'h0 : _GEN_637; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_639 = 10'h27f == io_inputs_0 ? 7'h0 : _GEN_638; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_640 = 10'h280 == io_inputs_0 ? 7'h0 : _GEN_639; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_641 = 10'h281 == io_inputs_0 ? 7'h0 : _GEN_640; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_642 = 10'h282 == io_inputs_0 ? 7'h0 : _GEN_641; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_643 = 10'h283 == io_inputs_0 ? 7'h0 : _GEN_642; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_644 = 10'h284 == io_inputs_0 ? 7'h0 : _GEN_643; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_645 = 10'h285 == io_inputs_0 ? 7'h0 : _GEN_644; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_646 = 10'h286 == io_inputs_0 ? 7'h0 : _GEN_645; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_647 = 10'h287 == io_inputs_0 ? 7'h0 : _GEN_646; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_648 = 10'h288 == io_inputs_0 ? 7'h0 : _GEN_647; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_649 = 10'h289 == io_inputs_0 ? 7'h0 : _GEN_648; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_650 = 10'h28a == io_inputs_0 ? 7'h0 : _GEN_649; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_651 = 10'h28b == io_inputs_0 ? 7'h0 : _GEN_650; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_652 = 10'h28c == io_inputs_0 ? 7'h0 : _GEN_651; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_653 = 10'h28d == io_inputs_0 ? 7'h0 : _GEN_652; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_654 = 10'h28e == io_inputs_0 ? 7'h0 : _GEN_653; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_655 = 10'h28f == io_inputs_0 ? 7'h0 : _GEN_654; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_656 = 10'h290 == io_inputs_0 ? 7'h0 : _GEN_655; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_657 = 10'h291 == io_inputs_0 ? 7'h0 : _GEN_656; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_658 = 10'h292 == io_inputs_0 ? 7'h0 : _GEN_657; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_659 = 10'h293 == io_inputs_0 ? 7'h0 : _GEN_658; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_660 = 10'h294 == io_inputs_0 ? 7'h0 : _GEN_659; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_661 = 10'h295 == io_inputs_0 ? 7'h0 : _GEN_660; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_662 = 10'h296 == io_inputs_0 ? 7'h0 : _GEN_661; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_663 = 10'h297 == io_inputs_0 ? 7'h0 : _GEN_662; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_664 = 10'h298 == io_inputs_0 ? 7'h0 : _GEN_663; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_665 = 10'h299 == io_inputs_0 ? 7'h0 : _GEN_664; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_666 = 10'h29a == io_inputs_0 ? 7'h0 : _GEN_665; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_667 = 10'h29b == io_inputs_0 ? 7'h0 : _GEN_666; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_668 = 10'h29c == io_inputs_0 ? 7'h0 : _GEN_667; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_669 = 10'h29d == io_inputs_0 ? 7'h0 : _GEN_668; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_670 = 10'h29e == io_inputs_0 ? 7'h0 : _GEN_669; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_671 = 10'h29f == io_inputs_0 ? 7'h0 : _GEN_670; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_672 = 10'h2a0 == io_inputs_0 ? 7'h0 : _GEN_671; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_673 = 10'h2a1 == io_inputs_0 ? 7'h0 : _GEN_672; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_674 = 10'h2a2 == io_inputs_0 ? 7'h0 : _GEN_673; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_675 = 10'h2a3 == io_inputs_0 ? 7'h0 : _GEN_674; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_676 = 10'h2a4 == io_inputs_0 ? 7'h0 : _GEN_675; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_677 = 10'h2a5 == io_inputs_0 ? 7'h0 : _GEN_676; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_678 = 10'h2a6 == io_inputs_0 ? 7'h0 : _GEN_677; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_679 = 10'h2a7 == io_inputs_0 ? 7'h0 : _GEN_678; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_680 = 10'h2a8 == io_inputs_0 ? 7'h0 : _GEN_679; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_681 = 10'h2a9 == io_inputs_0 ? 7'h0 : _GEN_680; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_682 = 10'h2aa == io_inputs_0 ? 7'h0 : _GEN_681; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_683 = 10'h2ab == io_inputs_0 ? 7'h0 : _GEN_682; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_684 = 10'h2ac == io_inputs_0 ? 7'h0 : _GEN_683; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_685 = 10'h2ad == io_inputs_0 ? 7'h0 : _GEN_684; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_686 = 10'h2ae == io_inputs_0 ? 7'h0 : _GEN_685; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_687 = 10'h2af == io_inputs_0 ? 7'h0 : _GEN_686; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_688 = 10'h2b0 == io_inputs_0 ? 7'h0 : _GEN_687; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_689 = 10'h2b1 == io_inputs_0 ? 7'h0 : _GEN_688; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_690 = 10'h2b2 == io_inputs_0 ? 7'h0 : _GEN_689; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_691 = 10'h2b3 == io_inputs_0 ? 7'h0 : _GEN_690; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_692 = 10'h2b4 == io_inputs_0 ? 7'h0 : _GEN_691; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_693 = 10'h2b5 == io_inputs_0 ? 7'h0 : _GEN_692; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_694 = 10'h2b6 == io_inputs_0 ? 7'h0 : _GEN_693; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_695 = 10'h2b7 == io_inputs_0 ? 7'h0 : _GEN_694; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_696 = 10'h2b8 == io_inputs_0 ? 7'h0 : _GEN_695; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_697 = 10'h2b9 == io_inputs_0 ? 7'h0 : _GEN_696; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_698 = 10'h2ba == io_inputs_0 ? 7'h0 : _GEN_697; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_699 = 10'h2bb == io_inputs_0 ? 7'h0 : _GEN_698; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_700 = 10'h2bc == io_inputs_0 ? 7'h0 : _GEN_699; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_701 = 10'h2bd == io_inputs_0 ? 7'h0 : _GEN_700; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_702 = 10'h2be == io_inputs_0 ? 7'h0 : _GEN_701; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_703 = 10'h2bf == io_inputs_0 ? 7'h0 : _GEN_702; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_704 = 10'h2c0 == io_inputs_0 ? 7'h0 : _GEN_703; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_705 = 10'h2c1 == io_inputs_0 ? 7'h0 : _GEN_704; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_706 = 10'h2c2 == io_inputs_0 ? 7'h0 : _GEN_705; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_707 = 10'h2c3 == io_inputs_0 ? 7'h0 : _GEN_706; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_708 = 10'h2c4 == io_inputs_0 ? 7'h0 : _GEN_707; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_709 = 10'h2c5 == io_inputs_0 ? 7'h0 : _GEN_708; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_710 = 10'h2c6 == io_inputs_0 ? 7'h0 : _GEN_709; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_711 = 10'h2c7 == io_inputs_0 ? 7'h0 : _GEN_710; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_712 = 10'h2c8 == io_inputs_0 ? 7'h0 : _GEN_711; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_713 = 10'h2c9 == io_inputs_0 ? 7'h0 : _GEN_712; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_714 = 10'h2ca == io_inputs_0 ? 7'h0 : _GEN_713; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_715 = 10'h2cb == io_inputs_0 ? 7'h0 : _GEN_714; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_716 = 10'h2cc == io_inputs_0 ? 7'h0 : _GEN_715; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_717 = 10'h2cd == io_inputs_0 ? 7'h0 : _GEN_716; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_718 = 10'h2ce == io_inputs_0 ? 7'h0 : _GEN_717; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_719 = 10'h2cf == io_inputs_0 ? 7'h0 : _GEN_718; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_720 = 10'h2d0 == io_inputs_0 ? 7'h0 : _GEN_719; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_721 = 10'h2d1 == io_inputs_0 ? 7'h0 : _GEN_720; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_722 = 10'h2d2 == io_inputs_0 ? 7'h0 : _GEN_721; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_723 = 10'h2d3 == io_inputs_0 ? 7'h0 : _GEN_722; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_724 = 10'h2d4 == io_inputs_0 ? 7'h0 : _GEN_723; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_725 = 10'h2d5 == io_inputs_0 ? 7'h0 : _GEN_724; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_726 = 10'h2d6 == io_inputs_0 ? 7'h0 : _GEN_725; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_727 = 10'h2d7 == io_inputs_0 ? 7'h0 : _GEN_726; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_728 = 10'h2d8 == io_inputs_0 ? 7'h0 : _GEN_727; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_729 = 10'h2d9 == io_inputs_0 ? 7'h0 : _GEN_728; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_730 = 10'h2da == io_inputs_0 ? 7'h0 : _GEN_729; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_731 = 10'h2db == io_inputs_0 ? 7'h0 : _GEN_730; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_732 = 10'h2dc == io_inputs_0 ? 7'h0 : _GEN_731; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_733 = 10'h2dd == io_inputs_0 ? 7'h0 : _GEN_732; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_734 = 10'h2de == io_inputs_0 ? 7'h0 : _GEN_733; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_735 = 10'h2df == io_inputs_0 ? 7'h0 : _GEN_734; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_736 = 10'h2e0 == io_inputs_0 ? 7'h0 : _GEN_735; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_737 = 10'h2e1 == io_inputs_0 ? 7'h0 : _GEN_736; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_738 = 10'h2e2 == io_inputs_0 ? 7'h0 : _GEN_737; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_739 = 10'h2e3 == io_inputs_0 ? 7'h0 : _GEN_738; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_740 = 10'h2e4 == io_inputs_0 ? 7'h0 : _GEN_739; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_741 = 10'h2e5 == io_inputs_0 ? 7'h0 : _GEN_740; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_742 = 10'h2e6 == io_inputs_0 ? 7'h0 : _GEN_741; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_743 = 10'h2e7 == io_inputs_0 ? 7'h0 : _GEN_742; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_744 = 10'h2e8 == io_inputs_0 ? 7'h0 : _GEN_743; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_745 = 10'h2e9 == io_inputs_0 ? 7'h0 : _GEN_744; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_746 = 10'h2ea == io_inputs_0 ? 7'h0 : _GEN_745; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_747 = 10'h2eb == io_inputs_0 ? 7'h0 : _GEN_746; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_748 = 10'h2ec == io_inputs_0 ? 7'h0 : _GEN_747; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_749 = 10'h2ed == io_inputs_0 ? 7'h0 : _GEN_748; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_750 = 10'h2ee == io_inputs_0 ? 7'h0 : _GEN_749; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_751 = 10'h2ef == io_inputs_0 ? 7'h0 : _GEN_750; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_752 = 10'h2f0 == io_inputs_0 ? 7'h0 : _GEN_751; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_753 = 10'h2f1 == io_inputs_0 ? 7'h0 : _GEN_752; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_754 = 10'h2f2 == io_inputs_0 ? 7'h0 : _GEN_753; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_755 = 10'h2f3 == io_inputs_0 ? 7'h0 : _GEN_754; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_756 = 10'h2f4 == io_inputs_0 ? 7'h0 : _GEN_755; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_757 = 10'h2f5 == io_inputs_0 ? 7'h0 : _GEN_756; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_758 = 10'h2f6 == io_inputs_0 ? 7'h0 : _GEN_757; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_759 = 10'h2f7 == io_inputs_0 ? 7'h0 : _GEN_758; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_760 = 10'h2f8 == io_inputs_0 ? 7'h0 : _GEN_759; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_761 = 10'h2f9 == io_inputs_0 ? 7'h0 : _GEN_760; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_762 = 10'h2fa == io_inputs_0 ? 7'h0 : _GEN_761; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_763 = 10'h2fb == io_inputs_0 ? 7'h0 : _GEN_762; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_764 = 10'h2fc == io_inputs_0 ? 7'h0 : _GEN_763; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_765 = 10'h2fd == io_inputs_0 ? 7'h0 : _GEN_764; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_766 = 10'h2fe == io_inputs_0 ? 7'h0 : _GEN_765; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_767 = 10'h2ff == io_inputs_0 ? 7'h0 : _GEN_766; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_768 = 10'h300 == io_inputs_0 ? 7'h0 : _GEN_767; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_769 = 10'h301 == io_inputs_0 ? 7'h0 : _GEN_768; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_770 = 10'h302 == io_inputs_0 ? 7'h0 : _GEN_769; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_771 = 10'h303 == io_inputs_0 ? 7'h0 : _GEN_770; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_772 = 10'h304 == io_inputs_0 ? 7'h0 : _GEN_771; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_773 = 10'h305 == io_inputs_0 ? 7'h0 : _GEN_772; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_774 = 10'h306 == io_inputs_0 ? 7'h0 : _GEN_773; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_775 = 10'h307 == io_inputs_0 ? 7'h0 : _GEN_774; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_776 = 10'h308 == io_inputs_0 ? 7'h0 : _GEN_775; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_777 = 10'h309 == io_inputs_0 ? 7'h0 : _GEN_776; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_778 = 10'h30a == io_inputs_0 ? 7'h0 : _GEN_777; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_779 = 10'h30b == io_inputs_0 ? 7'h0 : _GEN_778; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_780 = 10'h30c == io_inputs_0 ? 7'h0 : _GEN_779; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_781 = 10'h30d == io_inputs_0 ? 7'h0 : _GEN_780; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_782 = 10'h30e == io_inputs_0 ? 7'h0 : _GEN_781; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_783 = 10'h30f == io_inputs_0 ? 7'h0 : _GEN_782; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_784 = 10'h310 == io_inputs_0 ? 7'h0 : _GEN_783; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_785 = 10'h311 == io_inputs_0 ? 7'h0 : _GEN_784; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_786 = 10'h312 == io_inputs_0 ? 7'h0 : _GEN_785; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_787 = 10'h313 == io_inputs_0 ? 7'h0 : _GEN_786; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_788 = 10'h314 == io_inputs_0 ? 7'h0 : _GEN_787; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_789 = 10'h315 == io_inputs_0 ? 7'h0 : _GEN_788; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_790 = 10'h316 == io_inputs_0 ? 7'h0 : _GEN_789; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_791 = 10'h317 == io_inputs_0 ? 7'h0 : _GEN_790; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_792 = 10'h318 == io_inputs_0 ? 7'h0 : _GEN_791; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_793 = 10'h319 == io_inputs_0 ? 7'h0 : _GEN_792; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_794 = 10'h31a == io_inputs_0 ? 7'h0 : _GEN_793; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_795 = 10'h31b == io_inputs_0 ? 7'h0 : _GEN_794; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_796 = 10'h31c == io_inputs_0 ? 7'h0 : _GEN_795; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_797 = 10'h31d == io_inputs_0 ? 7'h0 : _GEN_796; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_798 = 10'h31e == io_inputs_0 ? 7'h0 : _GEN_797; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_799 = 10'h31f == io_inputs_0 ? 7'h0 : _GEN_798; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_800 = 10'h320 == io_inputs_0 ? 7'h0 : _GEN_799; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_801 = 10'h321 == io_inputs_0 ? 7'h0 : _GEN_800; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_802 = 10'h322 == io_inputs_0 ? 7'h0 : _GEN_801; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_803 = 10'h323 == io_inputs_0 ? 7'h0 : _GEN_802; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_804 = 10'h324 == io_inputs_0 ? 7'h0 : _GEN_803; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_805 = 10'h325 == io_inputs_0 ? 7'h0 : _GEN_804; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_806 = 10'h326 == io_inputs_0 ? 7'h0 : _GEN_805; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_807 = 10'h327 == io_inputs_0 ? 7'h0 : _GEN_806; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_808 = 10'h328 == io_inputs_0 ? 7'h0 : _GEN_807; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_809 = 10'h329 == io_inputs_0 ? 7'h0 : _GEN_808; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_810 = 10'h32a == io_inputs_0 ? 7'h0 : _GEN_809; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_811 = 10'h32b == io_inputs_0 ? 7'h0 : _GEN_810; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_812 = 10'h32c == io_inputs_0 ? 7'h0 : _GEN_811; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_813 = 10'h32d == io_inputs_0 ? 7'h0 : _GEN_812; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_814 = 10'h32e == io_inputs_0 ? 7'h0 : _GEN_813; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_815 = 10'h32f == io_inputs_0 ? 7'h0 : _GEN_814; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_816 = 10'h330 == io_inputs_0 ? 7'h0 : _GEN_815; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_817 = 10'h331 == io_inputs_0 ? 7'h0 : _GEN_816; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_818 = 10'h332 == io_inputs_0 ? 7'h0 : _GEN_817; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_819 = 10'h333 == io_inputs_0 ? 7'h0 : _GEN_818; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_820 = 10'h334 == io_inputs_0 ? 7'h0 : _GEN_819; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_821 = 10'h335 == io_inputs_0 ? 7'h0 : _GEN_820; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_822 = 10'h336 == io_inputs_0 ? 7'h0 : _GEN_821; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_823 = 10'h337 == io_inputs_0 ? 7'h0 : _GEN_822; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_824 = 10'h338 == io_inputs_0 ? 7'h0 : _GEN_823; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_825 = 10'h339 == io_inputs_0 ? 7'h0 : _GEN_824; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_826 = 10'h33a == io_inputs_0 ? 7'h0 : _GEN_825; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_827 = 10'h33b == io_inputs_0 ? 7'h0 : _GEN_826; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_828 = 10'h33c == io_inputs_0 ? 7'h0 : _GEN_827; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_829 = 10'h33d == io_inputs_0 ? 7'h0 : _GEN_828; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_830 = 10'h33e == io_inputs_0 ? 7'h0 : _GEN_829; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_831 = 10'h33f == io_inputs_0 ? 7'h0 : _GEN_830; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_832 = 10'h340 == io_inputs_0 ? 7'h0 : _GEN_831; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_833 = 10'h341 == io_inputs_0 ? 7'h0 : _GEN_832; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_834 = 10'h342 == io_inputs_0 ? 7'h0 : _GEN_833; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_835 = 10'h343 == io_inputs_0 ? 7'h0 : _GEN_834; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_836 = 10'h344 == io_inputs_0 ? 7'h0 : _GEN_835; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_837 = 10'h345 == io_inputs_0 ? 7'h0 : _GEN_836; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_838 = 10'h346 == io_inputs_0 ? 7'h0 : _GEN_837; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_839 = 10'h347 == io_inputs_0 ? 7'h0 : _GEN_838; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_840 = 10'h348 == io_inputs_0 ? 7'h0 : _GEN_839; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_841 = 10'h349 == io_inputs_0 ? 7'h0 : _GEN_840; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_842 = 10'h34a == io_inputs_0 ? 7'h0 : _GEN_841; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_843 = 10'h34b == io_inputs_0 ? 7'h0 : _GEN_842; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_844 = 10'h34c == io_inputs_0 ? 7'h0 : _GEN_843; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_845 = 10'h34d == io_inputs_0 ? 7'h0 : _GEN_844; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_846 = 10'h34e == io_inputs_0 ? 7'h0 : _GEN_845; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_847 = 10'h34f == io_inputs_0 ? 7'h0 : _GEN_846; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_848 = 10'h350 == io_inputs_0 ? 7'h0 : _GEN_847; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_849 = 10'h351 == io_inputs_0 ? 7'h0 : _GEN_848; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_850 = 10'h352 == io_inputs_0 ? 7'h0 : _GEN_849; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_851 = 10'h353 == io_inputs_0 ? 7'h0 : _GEN_850; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_852 = 10'h354 == io_inputs_0 ? 7'h0 : _GEN_851; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_853 = 10'h355 == io_inputs_0 ? 7'h0 : _GEN_852; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_854 = 10'h356 == io_inputs_0 ? 7'h0 : _GEN_853; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_855 = 10'h357 == io_inputs_0 ? 7'h0 : _GEN_854; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_856 = 10'h358 == io_inputs_0 ? 7'h0 : _GEN_855; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_857 = 10'h359 == io_inputs_0 ? 7'h0 : _GEN_856; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_858 = 10'h35a == io_inputs_0 ? 7'h0 : _GEN_857; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_859 = 10'h35b == io_inputs_0 ? 7'h0 : _GEN_858; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_860 = 10'h35c == io_inputs_0 ? 7'h0 : _GEN_859; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_861 = 10'h35d == io_inputs_0 ? 7'h0 : _GEN_860; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_862 = 10'h35e == io_inputs_0 ? 7'h0 : _GEN_861; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_863 = 10'h35f == io_inputs_0 ? 7'h0 : _GEN_862; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_864 = 10'h360 == io_inputs_0 ? 7'h0 : _GEN_863; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_865 = 10'h361 == io_inputs_0 ? 7'h0 : _GEN_864; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_866 = 10'h362 == io_inputs_0 ? 7'h0 : _GEN_865; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_867 = 10'h363 == io_inputs_0 ? 7'h0 : _GEN_866; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_868 = 10'h364 == io_inputs_0 ? 7'h0 : _GEN_867; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_869 = 10'h365 == io_inputs_0 ? 7'h0 : _GEN_868; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_870 = 10'h366 == io_inputs_0 ? 7'h0 : _GEN_869; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_871 = 10'h367 == io_inputs_0 ? 7'h0 : _GEN_870; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_872 = 10'h368 == io_inputs_0 ? 7'h0 : _GEN_871; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_873 = 10'h369 == io_inputs_0 ? 7'h0 : _GEN_872; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_874 = 10'h36a == io_inputs_0 ? 7'h0 : _GEN_873; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_875 = 10'h36b == io_inputs_0 ? 7'h0 : _GEN_874; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_876 = 10'h36c == io_inputs_0 ? 7'h0 : _GEN_875; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_877 = 10'h36d == io_inputs_0 ? 7'h0 : _GEN_876; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_878 = 10'h36e == io_inputs_0 ? 7'h0 : _GEN_877; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_879 = 10'h36f == io_inputs_0 ? 7'h0 : _GEN_878; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_880 = 10'h370 == io_inputs_0 ? 7'h0 : _GEN_879; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_881 = 10'h371 == io_inputs_0 ? 7'h0 : _GEN_880; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_882 = 10'h372 == io_inputs_0 ? 7'h0 : _GEN_881; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_883 = 10'h373 == io_inputs_0 ? 7'h0 : _GEN_882; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_884 = 10'h374 == io_inputs_0 ? 7'h0 : _GEN_883; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_885 = 10'h375 == io_inputs_0 ? 7'h0 : _GEN_884; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_886 = 10'h376 == io_inputs_0 ? 7'h0 : _GEN_885; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_887 = 10'h377 == io_inputs_0 ? 7'h0 : _GEN_886; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_888 = 10'h378 == io_inputs_0 ? 7'h0 : _GEN_887; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_889 = 10'h379 == io_inputs_0 ? 7'h0 : _GEN_888; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_890 = 10'h37a == io_inputs_0 ? 7'h0 : _GEN_889; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_891 = 10'h37b == io_inputs_0 ? 7'h0 : _GEN_890; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_892 = 10'h37c == io_inputs_0 ? 7'h0 : _GEN_891; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_893 = 10'h37d == io_inputs_0 ? 7'h0 : _GEN_892; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_894 = 10'h37e == io_inputs_0 ? 7'h0 : _GEN_893; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_895 = 10'h37f == io_inputs_0 ? 7'h0 : _GEN_894; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_896 = 10'h380 == io_inputs_0 ? 7'h0 : _GEN_895; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_897 = 10'h381 == io_inputs_0 ? 7'h0 : _GEN_896; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_898 = 10'h382 == io_inputs_0 ? 7'h0 : _GEN_897; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_899 = 10'h383 == io_inputs_0 ? 7'h0 : _GEN_898; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_900 = 10'h384 == io_inputs_0 ? 7'h0 : _GEN_899; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_901 = 10'h385 == io_inputs_0 ? 7'h0 : _GEN_900; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_902 = 10'h386 == io_inputs_0 ? 7'h0 : _GEN_901; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_903 = 10'h387 == io_inputs_0 ? 7'h0 : _GEN_902; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_904 = 10'h388 == io_inputs_0 ? 7'h0 : _GEN_903; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_905 = 10'h389 == io_inputs_0 ? 7'h0 : _GEN_904; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_906 = 10'h38a == io_inputs_0 ? 7'h0 : _GEN_905; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_907 = 10'h38b == io_inputs_0 ? 7'h0 : _GEN_906; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_908 = 10'h38c == io_inputs_0 ? 7'h0 : _GEN_907; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_909 = 10'h38d == io_inputs_0 ? 7'h0 : _GEN_908; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_910 = 10'h38e == io_inputs_0 ? 7'h0 : _GEN_909; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_911 = 10'h38f == io_inputs_0 ? 7'h0 : _GEN_910; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_912 = 10'h390 == io_inputs_0 ? 7'h0 : _GEN_911; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_913 = 10'h391 == io_inputs_0 ? 7'h0 : _GEN_912; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_914 = 10'h392 == io_inputs_0 ? 7'h0 : _GEN_913; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_915 = 10'h393 == io_inputs_0 ? 7'h0 : _GEN_914; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_916 = 10'h394 == io_inputs_0 ? 7'h0 : _GEN_915; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_917 = 10'h395 == io_inputs_0 ? 7'h0 : _GEN_916; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_918 = 10'h396 == io_inputs_0 ? 7'h0 : _GEN_917; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_919 = 10'h397 == io_inputs_0 ? 7'h0 : _GEN_918; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_920 = 10'h398 == io_inputs_0 ? 7'h0 : _GEN_919; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_921 = 10'h399 == io_inputs_0 ? 7'h0 : _GEN_920; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_922 = 10'h39a == io_inputs_0 ? 7'h0 : _GEN_921; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_923 = 10'h39b == io_inputs_0 ? 7'h0 : _GEN_922; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_924 = 10'h39c == io_inputs_0 ? 7'h0 : _GEN_923; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_925 = 10'h39d == io_inputs_0 ? 7'h0 : _GEN_924; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_926 = 10'h39e == io_inputs_0 ? 7'h0 : _GEN_925; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_927 = 10'h39f == io_inputs_0 ? 7'h0 : _GEN_926; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_928 = 10'h3a0 == io_inputs_0 ? 7'h0 : _GEN_927; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_929 = 10'h3a1 == io_inputs_0 ? 7'h0 : _GEN_928; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_930 = 10'h3a2 == io_inputs_0 ? 7'h0 : _GEN_929; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_931 = 10'h3a3 == io_inputs_0 ? 7'h0 : _GEN_930; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_932 = 10'h3a4 == io_inputs_0 ? 7'h0 : _GEN_931; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_933 = 10'h3a5 == io_inputs_0 ? 7'h0 : _GEN_932; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_934 = 10'h3a6 == io_inputs_0 ? 7'h0 : _GEN_933; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_935 = 10'h3a7 == io_inputs_0 ? 7'h0 : _GEN_934; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_936 = 10'h3a8 == io_inputs_0 ? 7'h0 : _GEN_935; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_937 = 10'h3a9 == io_inputs_0 ? 7'h0 : _GEN_936; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_938 = 10'h3aa == io_inputs_0 ? 7'h0 : _GEN_937; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_939 = 10'h3ab == io_inputs_0 ? 7'h0 : _GEN_938; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_940 = 10'h3ac == io_inputs_0 ? 7'h0 : _GEN_939; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_941 = 10'h3ad == io_inputs_0 ? 7'h0 : _GEN_940; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_942 = 10'h3ae == io_inputs_0 ? 7'h0 : _GEN_941; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_943 = 10'h3af == io_inputs_0 ? 7'h0 : _GEN_942; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_944 = 10'h3b0 == io_inputs_0 ? 7'h0 : _GEN_943; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_945 = 10'h3b1 == io_inputs_0 ? 7'h0 : _GEN_944; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_946 = 10'h3b2 == io_inputs_0 ? 7'h0 : _GEN_945; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_947 = 10'h3b3 == io_inputs_0 ? 7'h0 : _GEN_946; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_948 = 10'h3b4 == io_inputs_0 ? 7'h0 : _GEN_947; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_949 = 10'h3b5 == io_inputs_0 ? 7'h0 : _GEN_948; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_950 = 10'h3b6 == io_inputs_0 ? 7'h0 : _GEN_949; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_951 = 10'h3b7 == io_inputs_0 ? 7'h0 : _GEN_950; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_952 = 10'h3b8 == io_inputs_0 ? 7'h0 : _GEN_951; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_953 = 10'h3b9 == io_inputs_0 ? 7'h0 : _GEN_952; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_954 = 10'h3ba == io_inputs_0 ? 7'h0 : _GEN_953; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_955 = 10'h3bb == io_inputs_0 ? 7'h0 : _GEN_954; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_956 = 10'h3bc == io_inputs_0 ? 7'h0 : _GEN_955; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_957 = 10'h3bd == io_inputs_0 ? 7'h0 : _GEN_956; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_958 = 10'h3be == io_inputs_0 ? 7'h0 : _GEN_957; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_959 = 10'h3bf == io_inputs_0 ? 7'h0 : _GEN_958; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_960 = 10'h3c0 == io_inputs_0 ? 7'h0 : _GEN_959; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_961 = 10'h3c1 == io_inputs_0 ? 7'h0 : _GEN_960; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_962 = 10'h3c2 == io_inputs_0 ? 7'h0 : _GEN_961; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_963 = 10'h3c3 == io_inputs_0 ? 7'h0 : _GEN_962; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_964 = 10'h3c4 == io_inputs_0 ? 7'h0 : _GEN_963; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_965 = 10'h3c5 == io_inputs_0 ? 7'h0 : _GEN_964; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_966 = 10'h3c6 == io_inputs_0 ? 7'h0 : _GEN_965; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_967 = 10'h3c7 == io_inputs_0 ? 7'h0 : _GEN_966; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_968 = 10'h3c8 == io_inputs_0 ? 7'h0 : _GEN_967; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_969 = 10'h3c9 == io_inputs_0 ? 7'h0 : _GEN_968; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_970 = 10'h3ca == io_inputs_0 ? 7'h0 : _GEN_969; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_971 = 10'h3cb == io_inputs_0 ? 7'h0 : _GEN_970; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_972 = 10'h3cc == io_inputs_0 ? 7'h0 : _GEN_971; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_973 = 10'h3cd == io_inputs_0 ? 7'h0 : _GEN_972; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_974 = 10'h3ce == io_inputs_0 ? 7'h0 : _GEN_973; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_975 = 10'h3cf == io_inputs_0 ? 7'h0 : _GEN_974; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_976 = 10'h3d0 == io_inputs_0 ? 7'h0 : _GEN_975; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_977 = 10'h3d1 == io_inputs_0 ? 7'h0 : _GEN_976; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_978 = 10'h3d2 == io_inputs_0 ? 7'h0 : _GEN_977; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_979 = 10'h3d3 == io_inputs_0 ? 7'h0 : _GEN_978; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_980 = 10'h3d4 == io_inputs_0 ? 7'h0 : _GEN_979; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_981 = 10'h3d5 == io_inputs_0 ? 7'h0 : _GEN_980; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_982 = 10'h3d6 == io_inputs_0 ? 7'h0 : _GEN_981; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_983 = 10'h3d7 == io_inputs_0 ? 7'h0 : _GEN_982; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_984 = 10'h3d8 == io_inputs_0 ? 7'h0 : _GEN_983; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_985 = 10'h3d9 == io_inputs_0 ? 7'h0 : _GEN_984; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_986 = 10'h3da == io_inputs_0 ? 7'h0 : _GEN_985; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_987 = 10'h3db == io_inputs_0 ? 7'h0 : _GEN_986; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_988 = 10'h3dc == io_inputs_0 ? 7'h0 : _GEN_987; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_989 = 10'h3dd == io_inputs_0 ? 7'h0 : _GEN_988; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_990 = 10'h3de == io_inputs_0 ? 7'h0 : _GEN_989; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_991 = 10'h3df == io_inputs_0 ? 7'h0 : _GEN_990; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_992 = 10'h3e0 == io_inputs_0 ? 7'h0 : _GEN_991; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_993 = 10'h3e1 == io_inputs_0 ? 7'h0 : _GEN_992; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_994 = 10'h3e2 == io_inputs_0 ? 7'h0 : _GEN_993; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_995 = 10'h3e3 == io_inputs_0 ? 7'h0 : _GEN_994; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_996 = 10'h3e4 == io_inputs_0 ? 7'h0 : _GEN_995; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_997 = 10'h3e5 == io_inputs_0 ? 7'h0 : _GEN_996; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_998 = 10'h3e6 == io_inputs_0 ? 7'h0 : _GEN_997; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_999 = 10'h3e7 == io_inputs_0 ? 7'h0 : _GEN_998; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1000 = 10'h3e8 == io_inputs_0 ? 7'h0 : _GEN_999; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1001 = 10'h3e9 == io_inputs_0 ? 7'h0 : _GEN_1000; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1002 = 10'h3ea == io_inputs_0 ? 7'h0 : _GEN_1001; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1003 = 10'h3eb == io_inputs_0 ? 7'h0 : _GEN_1002; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1004 = 10'h3ec == io_inputs_0 ? 7'h0 : _GEN_1003; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1005 = 10'h3ed == io_inputs_0 ? 7'h0 : _GEN_1004; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1006 = 10'h3ee == io_inputs_0 ? 7'h0 : _GEN_1005; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1007 = 10'h3ef == io_inputs_0 ? 7'h0 : _GEN_1006; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1008 = 10'h3f0 == io_inputs_0 ? 7'h0 : _GEN_1007; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1009 = 10'h3f1 == io_inputs_0 ? 7'h0 : _GEN_1008; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1010 = 10'h3f2 == io_inputs_0 ? 7'h0 : _GEN_1009; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1011 = 10'h3f3 == io_inputs_0 ? 7'h0 : _GEN_1010; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1012 = 10'h3f4 == io_inputs_0 ? 7'h0 : _GEN_1011; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1013 = 10'h3f5 == io_inputs_0 ? 7'h0 : _GEN_1012; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1014 = 10'h3f6 == io_inputs_0 ? 7'h0 : _GEN_1013; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1015 = 10'h3f7 == io_inputs_0 ? 7'h0 : _GEN_1014; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1016 = 10'h3f8 == io_inputs_0 ? 7'h0 : _GEN_1015; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1017 = 10'h3f9 == io_inputs_0 ? 7'h0 : _GEN_1016; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1018 = 10'h3fa == io_inputs_0 ? 7'h0 : _GEN_1017; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1019 = 10'h3fb == io_inputs_0 ? 7'h0 : _GEN_1018; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1020 = 10'h3fc == io_inputs_0 ? 7'h0 : _GEN_1019; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1075 = 10'h33 == io_inputs_0 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1076 = 10'h34 == io_inputs_0 ? 7'h2 : _GEN_1075; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1077 = 10'h35 == io_inputs_0 ? 7'h3 : _GEN_1076; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1078 = 10'h36 == io_inputs_0 ? 7'h4 : _GEN_1077; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1079 = 10'h37 == io_inputs_0 ? 7'h5 : _GEN_1078; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1080 = 10'h38 == io_inputs_0 ? 7'h6 : _GEN_1079; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1081 = 10'h39 == io_inputs_0 ? 7'h7 : _GEN_1080; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1082 = 10'h3a == io_inputs_0 ? 7'h8 : _GEN_1081; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1083 = 10'h3b == io_inputs_0 ? 7'h9 : _GEN_1082; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1084 = 10'h3c == io_inputs_0 ? 7'ha : _GEN_1083; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1085 = 10'h3d == io_inputs_0 ? 7'hb : _GEN_1084; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1086 = 10'h3e == io_inputs_0 ? 7'hc : _GEN_1085; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1087 = 10'h3f == io_inputs_0 ? 7'hd : _GEN_1086; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1088 = 10'h40 == io_inputs_0 ? 7'he : _GEN_1087; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1089 = 10'h41 == io_inputs_0 ? 7'hf : _GEN_1088; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1090 = 10'h42 == io_inputs_0 ? 7'h10 : _GEN_1089; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1091 = 10'h43 == io_inputs_0 ? 7'h11 : _GEN_1090; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1092 = 10'h44 == io_inputs_0 ? 7'h12 : _GEN_1091; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1093 = 10'h45 == io_inputs_0 ? 7'h13 : _GEN_1092; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1094 = 10'h46 == io_inputs_0 ? 7'h14 : _GEN_1093; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1095 = 10'h47 == io_inputs_0 ? 7'h15 : _GEN_1094; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1096 = 10'h48 == io_inputs_0 ? 7'h16 : _GEN_1095; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1097 = 10'h49 == io_inputs_0 ? 7'h17 : _GEN_1096; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1098 = 10'h4a == io_inputs_0 ? 7'h18 : _GEN_1097; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1099 = 10'h4b == io_inputs_0 ? 7'h19 : _GEN_1098; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1100 = 10'h4c == io_inputs_0 ? 7'h1a : _GEN_1099; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1101 = 10'h4d == io_inputs_0 ? 7'h1b : _GEN_1100; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1102 = 10'h4e == io_inputs_0 ? 7'h1c : _GEN_1101; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1103 = 10'h4f == io_inputs_0 ? 7'h1d : _GEN_1102; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1104 = 10'h50 == io_inputs_0 ? 7'h1e : _GEN_1103; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1105 = 10'h51 == io_inputs_0 ? 7'h1f : _GEN_1104; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1106 = 10'h52 == io_inputs_0 ? 7'h20 : _GEN_1105; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1107 = 10'h53 == io_inputs_0 ? 7'h21 : _GEN_1106; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1108 = 10'h54 == io_inputs_0 ? 7'h22 : _GEN_1107; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1109 = 10'h55 == io_inputs_0 ? 7'h23 : _GEN_1108; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1110 = 10'h56 == io_inputs_0 ? 7'h24 : _GEN_1109; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1111 = 10'h57 == io_inputs_0 ? 7'h25 : _GEN_1110; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1112 = 10'h58 == io_inputs_0 ? 7'h26 : _GEN_1111; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1113 = 10'h59 == io_inputs_0 ? 7'h27 : _GEN_1112; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1114 = 10'h5a == io_inputs_0 ? 7'h28 : _GEN_1113; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1115 = 10'h5b == io_inputs_0 ? 7'h29 : _GEN_1114; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1116 = 10'h5c == io_inputs_0 ? 7'h2a : _GEN_1115; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1117 = 10'h5d == io_inputs_0 ? 7'h2b : _GEN_1116; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1118 = 10'h5e == io_inputs_0 ? 7'h2c : _GEN_1117; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1119 = 10'h5f == io_inputs_0 ? 7'h2d : _GEN_1118; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1120 = 10'h60 == io_inputs_0 ? 7'h2e : _GEN_1119; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1121 = 10'h61 == io_inputs_0 ? 7'h2f : _GEN_1120; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1122 = 10'h62 == io_inputs_0 ? 7'h30 : _GEN_1121; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1123 = 10'h63 == io_inputs_0 ? 7'h31 : _GEN_1122; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1124 = 10'h64 == io_inputs_0 ? 7'h32 : _GEN_1123; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1125 = 10'h65 == io_inputs_0 ? 7'h33 : _GEN_1124; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1126 = 10'h66 == io_inputs_0 ? 7'h34 : _GEN_1125; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1127 = 10'h67 == io_inputs_0 ? 7'h35 : _GEN_1126; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1128 = 10'h68 == io_inputs_0 ? 7'h36 : _GEN_1127; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1129 = 10'h69 == io_inputs_0 ? 7'h37 : _GEN_1128; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1130 = 10'h6a == io_inputs_0 ? 7'h38 : _GEN_1129; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1131 = 10'h6b == io_inputs_0 ? 7'h39 : _GEN_1130; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1132 = 10'h6c == io_inputs_0 ? 7'h3a : _GEN_1131; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1133 = 10'h6d == io_inputs_0 ? 7'h3b : _GEN_1132; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1134 = 10'h6e == io_inputs_0 ? 7'h3c : _GEN_1133; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1135 = 10'h6f == io_inputs_0 ? 7'h3d : _GEN_1134; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1136 = 10'h70 == io_inputs_0 ? 7'h3e : _GEN_1135; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1137 = 10'h71 == io_inputs_0 ? 7'h3f : _GEN_1136; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1138 = 10'h72 == io_inputs_0 ? 7'h40 : _GEN_1137; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1139 = 10'h73 == io_inputs_0 ? 7'h41 : _GEN_1138; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1140 = 10'h74 == io_inputs_0 ? 7'h42 : _GEN_1139; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1141 = 10'h75 == io_inputs_0 ? 7'h43 : _GEN_1140; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1142 = 10'h76 == io_inputs_0 ? 7'h44 : _GEN_1141; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1143 = 10'h77 == io_inputs_0 ? 7'h45 : _GEN_1142; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1144 = 10'h78 == io_inputs_0 ? 7'h46 : _GEN_1143; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1145 = 10'h79 == io_inputs_0 ? 7'h47 : _GEN_1144; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1146 = 10'h7a == io_inputs_0 ? 7'h48 : _GEN_1145; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1147 = 10'h7b == io_inputs_0 ? 7'h49 : _GEN_1146; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1148 = 10'h7c == io_inputs_0 ? 7'h4a : _GEN_1147; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1149 = 10'h7d == io_inputs_0 ? 7'h4b : _GEN_1148; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1150 = 10'h7e == io_inputs_0 ? 7'h4c : _GEN_1149; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1151 = 10'h7f == io_inputs_0 ? 7'h4d : _GEN_1150; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1152 = 10'h80 == io_inputs_0 ? 7'h4e : _GEN_1151; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1153 = 10'h81 == io_inputs_0 ? 7'h4f : _GEN_1152; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1154 = 10'h82 == io_inputs_0 ? 7'h50 : _GEN_1153; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1155 = 10'h83 == io_inputs_0 ? 7'h51 : _GEN_1154; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1156 = 10'h84 == io_inputs_0 ? 7'h52 : _GEN_1155; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1157 = 10'h85 == io_inputs_0 ? 7'h53 : _GEN_1156; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1158 = 10'h86 == io_inputs_0 ? 7'h54 : _GEN_1157; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1159 = 10'h87 == io_inputs_0 ? 7'h55 : _GEN_1158; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1160 = 10'h88 == io_inputs_0 ? 7'h56 : _GEN_1159; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1161 = 10'h89 == io_inputs_0 ? 7'h57 : _GEN_1160; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1162 = 10'h8a == io_inputs_0 ? 7'h58 : _GEN_1161; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1163 = 10'h8b == io_inputs_0 ? 7'h59 : _GEN_1162; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1164 = 10'h8c == io_inputs_0 ? 7'h5a : _GEN_1163; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1165 = 10'h8d == io_inputs_0 ? 7'h5b : _GEN_1164; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1166 = 10'h8e == io_inputs_0 ? 7'h5c : _GEN_1165; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1167 = 10'h8f == io_inputs_0 ? 7'h5d : _GEN_1166; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1168 = 10'h90 == io_inputs_0 ? 7'h5e : _GEN_1167; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1169 = 10'h91 == io_inputs_0 ? 7'h5f : _GEN_1168; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1170 = 10'h92 == io_inputs_0 ? 7'h60 : _GEN_1169; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1171 = 10'h93 == io_inputs_0 ? 7'h61 : _GEN_1170; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1172 = 10'h94 == io_inputs_0 ? 7'h62 : _GEN_1171; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1173 = 10'h95 == io_inputs_0 ? 7'h63 : _GEN_1172; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1174 = 10'h96 == io_inputs_0 ? 7'h64 : _GEN_1173; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1175 = 10'h97 == io_inputs_0 ? 7'h64 : _GEN_1174; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1176 = 10'h98 == io_inputs_0 ? 7'h64 : _GEN_1175; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1177 = 10'h99 == io_inputs_0 ? 7'h64 : _GEN_1176; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1178 = 10'h9a == io_inputs_0 ? 7'h64 : _GEN_1177; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1179 = 10'h9b == io_inputs_0 ? 7'h64 : _GEN_1178; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1180 = 10'h9c == io_inputs_0 ? 7'h64 : _GEN_1179; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1181 = 10'h9d == io_inputs_0 ? 7'h64 : _GEN_1180; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1182 = 10'h9e == io_inputs_0 ? 7'h64 : _GEN_1181; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1183 = 10'h9f == io_inputs_0 ? 7'h64 : _GEN_1182; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1184 = 10'ha0 == io_inputs_0 ? 7'h64 : _GEN_1183; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1185 = 10'ha1 == io_inputs_0 ? 7'h64 : _GEN_1184; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1186 = 10'ha2 == io_inputs_0 ? 7'h64 : _GEN_1185; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1187 = 10'ha3 == io_inputs_0 ? 7'h64 : _GEN_1186; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1188 = 10'ha4 == io_inputs_0 ? 7'h64 : _GEN_1187; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1189 = 10'ha5 == io_inputs_0 ? 7'h64 : _GEN_1188; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1190 = 10'ha6 == io_inputs_0 ? 7'h64 : _GEN_1189; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1191 = 10'ha7 == io_inputs_0 ? 7'h64 : _GEN_1190; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1192 = 10'ha8 == io_inputs_0 ? 7'h64 : _GEN_1191; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1193 = 10'ha9 == io_inputs_0 ? 7'h64 : _GEN_1192; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1194 = 10'haa == io_inputs_0 ? 7'h64 : _GEN_1193; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1195 = 10'hab == io_inputs_0 ? 7'h64 : _GEN_1194; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1196 = 10'hac == io_inputs_0 ? 7'h64 : _GEN_1195; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1197 = 10'had == io_inputs_0 ? 7'h64 : _GEN_1196; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1198 = 10'hae == io_inputs_0 ? 7'h64 : _GEN_1197; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1199 = 10'haf == io_inputs_0 ? 7'h64 : _GEN_1198; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1200 = 10'hb0 == io_inputs_0 ? 7'h64 : _GEN_1199; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1201 = 10'hb1 == io_inputs_0 ? 7'h64 : _GEN_1200; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1202 = 10'hb2 == io_inputs_0 ? 7'h64 : _GEN_1201; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1203 = 10'hb3 == io_inputs_0 ? 7'h64 : _GEN_1202; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1204 = 10'hb4 == io_inputs_0 ? 7'h64 : _GEN_1203; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1205 = 10'hb5 == io_inputs_0 ? 7'h64 : _GEN_1204; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1206 = 10'hb6 == io_inputs_0 ? 7'h64 : _GEN_1205; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1207 = 10'hb7 == io_inputs_0 ? 7'h64 : _GEN_1206; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1208 = 10'hb8 == io_inputs_0 ? 7'h64 : _GEN_1207; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1209 = 10'hb9 == io_inputs_0 ? 7'h64 : _GEN_1208; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1210 = 10'hba == io_inputs_0 ? 7'h64 : _GEN_1209; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1211 = 10'hbb == io_inputs_0 ? 7'h64 : _GEN_1210; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1212 = 10'hbc == io_inputs_0 ? 7'h64 : _GEN_1211; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1213 = 10'hbd == io_inputs_0 ? 7'h64 : _GEN_1212; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1214 = 10'hbe == io_inputs_0 ? 7'h64 : _GEN_1213; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1215 = 10'hbf == io_inputs_0 ? 7'h64 : _GEN_1214; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1216 = 10'hc0 == io_inputs_0 ? 7'h64 : _GEN_1215; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1217 = 10'hc1 == io_inputs_0 ? 7'h64 : _GEN_1216; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1218 = 10'hc2 == io_inputs_0 ? 7'h64 : _GEN_1217; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1219 = 10'hc3 == io_inputs_0 ? 7'h64 : _GEN_1218; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1220 = 10'hc4 == io_inputs_0 ? 7'h64 : _GEN_1219; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1221 = 10'hc5 == io_inputs_0 ? 7'h64 : _GEN_1220; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1222 = 10'hc6 == io_inputs_0 ? 7'h64 : _GEN_1221; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1223 = 10'hc7 == io_inputs_0 ? 7'h64 : _GEN_1222; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1224 = 10'hc8 == io_inputs_0 ? 7'h64 : _GEN_1223; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1225 = 10'hc9 == io_inputs_0 ? 7'h63 : _GEN_1224; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1226 = 10'hca == io_inputs_0 ? 7'h62 : _GEN_1225; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1227 = 10'hcb == io_inputs_0 ? 7'h61 : _GEN_1226; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1228 = 10'hcc == io_inputs_0 ? 7'h60 : _GEN_1227; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1229 = 10'hcd == io_inputs_0 ? 7'h5f : _GEN_1228; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1230 = 10'hce == io_inputs_0 ? 7'h5e : _GEN_1229; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1231 = 10'hcf == io_inputs_0 ? 7'h5d : _GEN_1230; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1232 = 10'hd0 == io_inputs_0 ? 7'h5c : _GEN_1231; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1233 = 10'hd1 == io_inputs_0 ? 7'h5b : _GEN_1232; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1234 = 10'hd2 == io_inputs_0 ? 7'h5a : _GEN_1233; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1235 = 10'hd3 == io_inputs_0 ? 7'h59 : _GEN_1234; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1236 = 10'hd4 == io_inputs_0 ? 7'h58 : _GEN_1235; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1237 = 10'hd5 == io_inputs_0 ? 7'h57 : _GEN_1236; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1238 = 10'hd6 == io_inputs_0 ? 7'h56 : _GEN_1237; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1239 = 10'hd7 == io_inputs_0 ? 7'h55 : _GEN_1238; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1240 = 10'hd8 == io_inputs_0 ? 7'h54 : _GEN_1239; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1241 = 10'hd9 == io_inputs_0 ? 7'h53 : _GEN_1240; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1242 = 10'hda == io_inputs_0 ? 7'h52 : _GEN_1241; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1243 = 10'hdb == io_inputs_0 ? 7'h51 : _GEN_1242; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1244 = 10'hdc == io_inputs_0 ? 7'h50 : _GEN_1243; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1245 = 10'hdd == io_inputs_0 ? 7'h4f : _GEN_1244; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1246 = 10'hde == io_inputs_0 ? 7'h4e : _GEN_1245; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1247 = 10'hdf == io_inputs_0 ? 7'h4d : _GEN_1246; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1248 = 10'he0 == io_inputs_0 ? 7'h4c : _GEN_1247; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1249 = 10'he1 == io_inputs_0 ? 7'h4b : _GEN_1248; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1250 = 10'he2 == io_inputs_0 ? 7'h4a : _GEN_1249; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1251 = 10'he3 == io_inputs_0 ? 7'h49 : _GEN_1250; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1252 = 10'he4 == io_inputs_0 ? 7'h48 : _GEN_1251; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1253 = 10'he5 == io_inputs_0 ? 7'h47 : _GEN_1252; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1254 = 10'he6 == io_inputs_0 ? 7'h46 : _GEN_1253; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1255 = 10'he7 == io_inputs_0 ? 7'h45 : _GEN_1254; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1256 = 10'he8 == io_inputs_0 ? 7'h44 : _GEN_1255; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1257 = 10'he9 == io_inputs_0 ? 7'h43 : _GEN_1256; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1258 = 10'hea == io_inputs_0 ? 7'h42 : _GEN_1257; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1259 = 10'heb == io_inputs_0 ? 7'h41 : _GEN_1258; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1260 = 10'hec == io_inputs_0 ? 7'h40 : _GEN_1259; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1261 = 10'hed == io_inputs_0 ? 7'h3f : _GEN_1260; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1262 = 10'hee == io_inputs_0 ? 7'h3e : _GEN_1261; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1263 = 10'hef == io_inputs_0 ? 7'h3d : _GEN_1262; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1264 = 10'hf0 == io_inputs_0 ? 7'h3c : _GEN_1263; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1265 = 10'hf1 == io_inputs_0 ? 7'h3b : _GEN_1264; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1266 = 10'hf2 == io_inputs_0 ? 7'h3a : _GEN_1265; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1267 = 10'hf3 == io_inputs_0 ? 7'h39 : _GEN_1266; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1268 = 10'hf4 == io_inputs_0 ? 7'h38 : _GEN_1267; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1269 = 10'hf5 == io_inputs_0 ? 7'h37 : _GEN_1268; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1270 = 10'hf6 == io_inputs_0 ? 7'h36 : _GEN_1269; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1271 = 10'hf7 == io_inputs_0 ? 7'h35 : _GEN_1270; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1272 = 10'hf8 == io_inputs_0 ? 7'h34 : _GEN_1271; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1273 = 10'hf9 == io_inputs_0 ? 7'h33 : _GEN_1272; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1274 = 10'hfa == io_inputs_0 ? 7'h32 : _GEN_1273; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1275 = 10'hfb == io_inputs_0 ? 7'h31 : _GEN_1274; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1276 = 10'hfc == io_inputs_0 ? 7'h30 : _GEN_1275; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1277 = 10'hfd == io_inputs_0 ? 7'h2f : _GEN_1276; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1278 = 10'hfe == io_inputs_0 ? 7'h2e : _GEN_1277; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1279 = 10'hff == io_inputs_0 ? 7'h2d : _GEN_1278; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1280 = 10'h100 == io_inputs_0 ? 7'h2c : _GEN_1279; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1281 = 10'h101 == io_inputs_0 ? 7'h2b : _GEN_1280; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1282 = 10'h102 == io_inputs_0 ? 7'h2a : _GEN_1281; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1283 = 10'h103 == io_inputs_0 ? 7'h29 : _GEN_1282; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1284 = 10'h104 == io_inputs_0 ? 7'h28 : _GEN_1283; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1285 = 10'h105 == io_inputs_0 ? 7'h27 : _GEN_1284; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1286 = 10'h106 == io_inputs_0 ? 7'h26 : _GEN_1285; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1287 = 10'h107 == io_inputs_0 ? 7'h25 : _GEN_1286; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1288 = 10'h108 == io_inputs_0 ? 7'h24 : _GEN_1287; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1289 = 10'h109 == io_inputs_0 ? 7'h23 : _GEN_1288; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1290 = 10'h10a == io_inputs_0 ? 7'h22 : _GEN_1289; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1291 = 10'h10b == io_inputs_0 ? 7'h21 : _GEN_1290; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1292 = 10'h10c == io_inputs_0 ? 7'h20 : _GEN_1291; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1293 = 10'h10d == io_inputs_0 ? 7'h1f : _GEN_1292; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1294 = 10'h10e == io_inputs_0 ? 7'h1e : _GEN_1293; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1295 = 10'h10f == io_inputs_0 ? 7'h1d : _GEN_1294; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1296 = 10'h110 == io_inputs_0 ? 7'h1c : _GEN_1295; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1297 = 10'h111 == io_inputs_0 ? 7'h1b : _GEN_1296; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1298 = 10'h112 == io_inputs_0 ? 7'h1a : _GEN_1297; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1299 = 10'h113 == io_inputs_0 ? 7'h19 : _GEN_1298; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1300 = 10'h114 == io_inputs_0 ? 7'h18 : _GEN_1299; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1301 = 10'h115 == io_inputs_0 ? 7'h17 : _GEN_1300; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1302 = 10'h116 == io_inputs_0 ? 7'h16 : _GEN_1301; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1303 = 10'h117 == io_inputs_0 ? 7'h15 : _GEN_1302; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1304 = 10'h118 == io_inputs_0 ? 7'h14 : _GEN_1303; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1305 = 10'h119 == io_inputs_0 ? 7'h13 : _GEN_1304; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1306 = 10'h11a == io_inputs_0 ? 7'h12 : _GEN_1305; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1307 = 10'h11b == io_inputs_0 ? 7'h11 : _GEN_1306; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1308 = 10'h11c == io_inputs_0 ? 7'h10 : _GEN_1307; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1309 = 10'h11d == io_inputs_0 ? 7'hf : _GEN_1308; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1310 = 10'h11e == io_inputs_0 ? 7'he : _GEN_1309; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1311 = 10'h11f == io_inputs_0 ? 7'hd : _GEN_1310; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1312 = 10'h120 == io_inputs_0 ? 7'hc : _GEN_1311; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1313 = 10'h121 == io_inputs_0 ? 7'hb : _GEN_1312; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1314 = 10'h122 == io_inputs_0 ? 7'ha : _GEN_1313; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1315 = 10'h123 == io_inputs_0 ? 7'h9 : _GEN_1314; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1316 = 10'h124 == io_inputs_0 ? 7'h8 : _GEN_1315; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1317 = 10'h125 == io_inputs_0 ? 7'h7 : _GEN_1316; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1318 = 10'h126 == io_inputs_0 ? 7'h6 : _GEN_1317; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1319 = 10'h127 == io_inputs_0 ? 7'h5 : _GEN_1318; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1320 = 10'h128 == io_inputs_0 ? 7'h4 : _GEN_1319; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1321 = 10'h129 == io_inputs_0 ? 7'h3 : _GEN_1320; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1322 = 10'h12a == io_inputs_0 ? 7'h2 : _GEN_1321; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1323 = 10'h12b == io_inputs_0 ? 7'h1 : _GEN_1322; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1324 = 10'h12c == io_inputs_0 ? 7'h0 : _GEN_1323; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1325 = 10'h12d == io_inputs_0 ? 7'h0 : _GEN_1324; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1326 = 10'h12e == io_inputs_0 ? 7'h0 : _GEN_1325; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1327 = 10'h12f == io_inputs_0 ? 7'h0 : _GEN_1326; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1328 = 10'h130 == io_inputs_0 ? 7'h0 : _GEN_1327; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1329 = 10'h131 == io_inputs_0 ? 7'h0 : _GEN_1328; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1330 = 10'h132 == io_inputs_0 ? 7'h0 : _GEN_1329; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1331 = 10'h133 == io_inputs_0 ? 7'h0 : _GEN_1330; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1332 = 10'h134 == io_inputs_0 ? 7'h0 : _GEN_1331; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1333 = 10'h135 == io_inputs_0 ? 7'h0 : _GEN_1332; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1334 = 10'h136 == io_inputs_0 ? 7'h0 : _GEN_1333; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1335 = 10'h137 == io_inputs_0 ? 7'h0 : _GEN_1334; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1336 = 10'h138 == io_inputs_0 ? 7'h0 : _GEN_1335; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1337 = 10'h139 == io_inputs_0 ? 7'h0 : _GEN_1336; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1338 = 10'h13a == io_inputs_0 ? 7'h0 : _GEN_1337; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1339 = 10'h13b == io_inputs_0 ? 7'h0 : _GEN_1338; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1340 = 10'h13c == io_inputs_0 ? 7'h0 : _GEN_1339; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1341 = 10'h13d == io_inputs_0 ? 7'h0 : _GEN_1340; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1342 = 10'h13e == io_inputs_0 ? 7'h0 : _GEN_1341; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1343 = 10'h13f == io_inputs_0 ? 7'h0 : _GEN_1342; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1344 = 10'h140 == io_inputs_0 ? 7'h0 : _GEN_1343; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1345 = 10'h141 == io_inputs_0 ? 7'h0 : _GEN_1344; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1346 = 10'h142 == io_inputs_0 ? 7'h0 : _GEN_1345; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1347 = 10'h143 == io_inputs_0 ? 7'h0 : _GEN_1346; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1348 = 10'h144 == io_inputs_0 ? 7'h0 : _GEN_1347; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1349 = 10'h145 == io_inputs_0 ? 7'h0 : _GEN_1348; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1350 = 10'h146 == io_inputs_0 ? 7'h0 : _GEN_1349; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1351 = 10'h147 == io_inputs_0 ? 7'h0 : _GEN_1350; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1352 = 10'h148 == io_inputs_0 ? 7'h0 : _GEN_1351; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1353 = 10'h149 == io_inputs_0 ? 7'h0 : _GEN_1352; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1354 = 10'h14a == io_inputs_0 ? 7'h0 : _GEN_1353; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1355 = 10'h14b == io_inputs_0 ? 7'h0 : _GEN_1354; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1356 = 10'h14c == io_inputs_0 ? 7'h0 : _GEN_1355; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1357 = 10'h14d == io_inputs_0 ? 7'h0 : _GEN_1356; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1358 = 10'h14e == io_inputs_0 ? 7'h0 : _GEN_1357; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1359 = 10'h14f == io_inputs_0 ? 7'h0 : _GEN_1358; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1360 = 10'h150 == io_inputs_0 ? 7'h0 : _GEN_1359; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1361 = 10'h151 == io_inputs_0 ? 7'h0 : _GEN_1360; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1362 = 10'h152 == io_inputs_0 ? 7'h0 : _GEN_1361; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1363 = 10'h153 == io_inputs_0 ? 7'h0 : _GEN_1362; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1364 = 10'h154 == io_inputs_0 ? 7'h0 : _GEN_1363; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1365 = 10'h155 == io_inputs_0 ? 7'h0 : _GEN_1364; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1366 = 10'h156 == io_inputs_0 ? 7'h0 : _GEN_1365; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1367 = 10'h157 == io_inputs_0 ? 7'h0 : _GEN_1366; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1368 = 10'h158 == io_inputs_0 ? 7'h0 : _GEN_1367; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1369 = 10'h159 == io_inputs_0 ? 7'h0 : _GEN_1368; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1370 = 10'h15a == io_inputs_0 ? 7'h0 : _GEN_1369; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1371 = 10'h15b == io_inputs_0 ? 7'h0 : _GEN_1370; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1372 = 10'h15c == io_inputs_0 ? 7'h0 : _GEN_1371; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1373 = 10'h15d == io_inputs_0 ? 7'h0 : _GEN_1372; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1374 = 10'h15e == io_inputs_0 ? 7'h0 : _GEN_1373; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1375 = 10'h15f == io_inputs_0 ? 7'h0 : _GEN_1374; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1376 = 10'h160 == io_inputs_0 ? 7'h0 : _GEN_1375; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1377 = 10'h161 == io_inputs_0 ? 7'h0 : _GEN_1376; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1378 = 10'h162 == io_inputs_0 ? 7'h0 : _GEN_1377; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1379 = 10'h163 == io_inputs_0 ? 7'h0 : _GEN_1378; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1380 = 10'h164 == io_inputs_0 ? 7'h0 : _GEN_1379; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1381 = 10'h165 == io_inputs_0 ? 7'h0 : _GEN_1380; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1382 = 10'h166 == io_inputs_0 ? 7'h0 : _GEN_1381; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1383 = 10'h167 == io_inputs_0 ? 7'h0 : _GEN_1382; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1384 = 10'h168 == io_inputs_0 ? 7'h0 : _GEN_1383; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1385 = 10'h169 == io_inputs_0 ? 7'h0 : _GEN_1384; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1386 = 10'h16a == io_inputs_0 ? 7'h0 : _GEN_1385; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1387 = 10'h16b == io_inputs_0 ? 7'h0 : _GEN_1386; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1388 = 10'h16c == io_inputs_0 ? 7'h0 : _GEN_1387; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1389 = 10'h16d == io_inputs_0 ? 7'h0 : _GEN_1388; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1390 = 10'h16e == io_inputs_0 ? 7'h0 : _GEN_1389; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1391 = 10'h16f == io_inputs_0 ? 7'h0 : _GEN_1390; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1392 = 10'h170 == io_inputs_0 ? 7'h0 : _GEN_1391; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1393 = 10'h171 == io_inputs_0 ? 7'h0 : _GEN_1392; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1394 = 10'h172 == io_inputs_0 ? 7'h0 : _GEN_1393; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1395 = 10'h173 == io_inputs_0 ? 7'h0 : _GEN_1394; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1396 = 10'h174 == io_inputs_0 ? 7'h0 : _GEN_1395; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1397 = 10'h175 == io_inputs_0 ? 7'h0 : _GEN_1396; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1398 = 10'h176 == io_inputs_0 ? 7'h0 : _GEN_1397; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1399 = 10'h177 == io_inputs_0 ? 7'h0 : _GEN_1398; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1400 = 10'h178 == io_inputs_0 ? 7'h0 : _GEN_1399; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1401 = 10'h179 == io_inputs_0 ? 7'h0 : _GEN_1400; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1402 = 10'h17a == io_inputs_0 ? 7'h0 : _GEN_1401; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1403 = 10'h17b == io_inputs_0 ? 7'h0 : _GEN_1402; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1404 = 10'h17c == io_inputs_0 ? 7'h0 : _GEN_1403; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1405 = 10'h17d == io_inputs_0 ? 7'h0 : _GEN_1404; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1406 = 10'h17e == io_inputs_0 ? 7'h0 : _GEN_1405; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1407 = 10'h17f == io_inputs_0 ? 7'h0 : _GEN_1406; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1408 = 10'h180 == io_inputs_0 ? 7'h0 : _GEN_1407; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1409 = 10'h181 == io_inputs_0 ? 7'h0 : _GEN_1408; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1410 = 10'h182 == io_inputs_0 ? 7'h0 : _GEN_1409; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1411 = 10'h183 == io_inputs_0 ? 7'h0 : _GEN_1410; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1412 = 10'h184 == io_inputs_0 ? 7'h0 : _GEN_1411; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1413 = 10'h185 == io_inputs_0 ? 7'h0 : _GEN_1412; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1414 = 10'h186 == io_inputs_0 ? 7'h0 : _GEN_1413; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1415 = 10'h187 == io_inputs_0 ? 7'h0 : _GEN_1414; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1416 = 10'h188 == io_inputs_0 ? 7'h0 : _GEN_1415; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1417 = 10'h189 == io_inputs_0 ? 7'h0 : _GEN_1416; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1418 = 10'h18a == io_inputs_0 ? 7'h0 : _GEN_1417; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1419 = 10'h18b == io_inputs_0 ? 7'h0 : _GEN_1418; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1420 = 10'h18c == io_inputs_0 ? 7'h0 : _GEN_1419; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1421 = 10'h18d == io_inputs_0 ? 7'h0 : _GEN_1420; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1422 = 10'h18e == io_inputs_0 ? 7'h0 : _GEN_1421; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1423 = 10'h18f == io_inputs_0 ? 7'h0 : _GEN_1422; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1424 = 10'h190 == io_inputs_0 ? 7'h0 : _GEN_1423; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1425 = 10'h191 == io_inputs_0 ? 7'h0 : _GEN_1424; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1426 = 10'h192 == io_inputs_0 ? 7'h0 : _GEN_1425; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1427 = 10'h193 == io_inputs_0 ? 7'h0 : _GEN_1426; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1428 = 10'h194 == io_inputs_0 ? 7'h0 : _GEN_1427; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1429 = 10'h195 == io_inputs_0 ? 7'h0 : _GEN_1428; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1430 = 10'h196 == io_inputs_0 ? 7'h0 : _GEN_1429; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1431 = 10'h197 == io_inputs_0 ? 7'h0 : _GEN_1430; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1432 = 10'h198 == io_inputs_0 ? 7'h0 : _GEN_1431; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1433 = 10'h199 == io_inputs_0 ? 7'h0 : _GEN_1432; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1434 = 10'h19a == io_inputs_0 ? 7'h0 : _GEN_1433; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1435 = 10'h19b == io_inputs_0 ? 7'h0 : _GEN_1434; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1436 = 10'h19c == io_inputs_0 ? 7'h0 : _GEN_1435; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1437 = 10'h19d == io_inputs_0 ? 7'h0 : _GEN_1436; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1438 = 10'h19e == io_inputs_0 ? 7'h0 : _GEN_1437; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1439 = 10'h19f == io_inputs_0 ? 7'h0 : _GEN_1438; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1440 = 10'h1a0 == io_inputs_0 ? 7'h0 : _GEN_1439; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1441 = 10'h1a1 == io_inputs_0 ? 7'h0 : _GEN_1440; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1442 = 10'h1a2 == io_inputs_0 ? 7'h0 : _GEN_1441; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1443 = 10'h1a3 == io_inputs_0 ? 7'h0 : _GEN_1442; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1444 = 10'h1a4 == io_inputs_0 ? 7'h0 : _GEN_1443; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1445 = 10'h1a5 == io_inputs_0 ? 7'h0 : _GEN_1444; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1446 = 10'h1a6 == io_inputs_0 ? 7'h0 : _GEN_1445; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1447 = 10'h1a7 == io_inputs_0 ? 7'h0 : _GEN_1446; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1448 = 10'h1a8 == io_inputs_0 ? 7'h0 : _GEN_1447; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1449 = 10'h1a9 == io_inputs_0 ? 7'h0 : _GEN_1448; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1450 = 10'h1aa == io_inputs_0 ? 7'h0 : _GEN_1449; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1451 = 10'h1ab == io_inputs_0 ? 7'h0 : _GEN_1450; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1452 = 10'h1ac == io_inputs_0 ? 7'h0 : _GEN_1451; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1453 = 10'h1ad == io_inputs_0 ? 7'h0 : _GEN_1452; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1454 = 10'h1ae == io_inputs_0 ? 7'h0 : _GEN_1453; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1455 = 10'h1af == io_inputs_0 ? 7'h0 : _GEN_1454; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1456 = 10'h1b0 == io_inputs_0 ? 7'h0 : _GEN_1455; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1457 = 10'h1b1 == io_inputs_0 ? 7'h0 : _GEN_1456; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1458 = 10'h1b2 == io_inputs_0 ? 7'h0 : _GEN_1457; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1459 = 10'h1b3 == io_inputs_0 ? 7'h0 : _GEN_1458; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1460 = 10'h1b4 == io_inputs_0 ? 7'h0 : _GEN_1459; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1461 = 10'h1b5 == io_inputs_0 ? 7'h0 : _GEN_1460; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1462 = 10'h1b6 == io_inputs_0 ? 7'h0 : _GEN_1461; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1463 = 10'h1b7 == io_inputs_0 ? 7'h0 : _GEN_1462; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1464 = 10'h1b8 == io_inputs_0 ? 7'h0 : _GEN_1463; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1465 = 10'h1b9 == io_inputs_0 ? 7'h0 : _GEN_1464; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1466 = 10'h1ba == io_inputs_0 ? 7'h0 : _GEN_1465; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1467 = 10'h1bb == io_inputs_0 ? 7'h0 : _GEN_1466; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1468 = 10'h1bc == io_inputs_0 ? 7'h0 : _GEN_1467; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1469 = 10'h1bd == io_inputs_0 ? 7'h0 : _GEN_1468; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1470 = 10'h1be == io_inputs_0 ? 7'h0 : _GEN_1469; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1471 = 10'h1bf == io_inputs_0 ? 7'h0 : _GEN_1470; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1472 = 10'h1c0 == io_inputs_0 ? 7'h0 : _GEN_1471; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1473 = 10'h1c1 == io_inputs_0 ? 7'h0 : _GEN_1472; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1474 = 10'h1c2 == io_inputs_0 ? 7'h0 : _GEN_1473; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1475 = 10'h1c3 == io_inputs_0 ? 7'h0 : _GEN_1474; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1476 = 10'h1c4 == io_inputs_0 ? 7'h0 : _GEN_1475; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1477 = 10'h1c5 == io_inputs_0 ? 7'h0 : _GEN_1476; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1478 = 10'h1c6 == io_inputs_0 ? 7'h0 : _GEN_1477; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1479 = 10'h1c7 == io_inputs_0 ? 7'h0 : _GEN_1478; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1480 = 10'h1c8 == io_inputs_0 ? 7'h0 : _GEN_1479; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1481 = 10'h1c9 == io_inputs_0 ? 7'h0 : _GEN_1480; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1482 = 10'h1ca == io_inputs_0 ? 7'h0 : _GEN_1481; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1483 = 10'h1cb == io_inputs_0 ? 7'h0 : _GEN_1482; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1484 = 10'h1cc == io_inputs_0 ? 7'h0 : _GEN_1483; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1485 = 10'h1cd == io_inputs_0 ? 7'h0 : _GEN_1484; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1486 = 10'h1ce == io_inputs_0 ? 7'h0 : _GEN_1485; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1487 = 10'h1cf == io_inputs_0 ? 7'h0 : _GEN_1486; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1488 = 10'h1d0 == io_inputs_0 ? 7'h0 : _GEN_1487; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1489 = 10'h1d1 == io_inputs_0 ? 7'h0 : _GEN_1488; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1490 = 10'h1d2 == io_inputs_0 ? 7'h0 : _GEN_1489; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1491 = 10'h1d3 == io_inputs_0 ? 7'h0 : _GEN_1490; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1492 = 10'h1d4 == io_inputs_0 ? 7'h0 : _GEN_1491; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1493 = 10'h1d5 == io_inputs_0 ? 7'h0 : _GEN_1492; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1494 = 10'h1d6 == io_inputs_0 ? 7'h0 : _GEN_1493; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1495 = 10'h1d7 == io_inputs_0 ? 7'h0 : _GEN_1494; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1496 = 10'h1d8 == io_inputs_0 ? 7'h0 : _GEN_1495; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1497 = 10'h1d9 == io_inputs_0 ? 7'h0 : _GEN_1496; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1498 = 10'h1da == io_inputs_0 ? 7'h0 : _GEN_1497; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1499 = 10'h1db == io_inputs_0 ? 7'h0 : _GEN_1498; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1500 = 10'h1dc == io_inputs_0 ? 7'h0 : _GEN_1499; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1501 = 10'h1dd == io_inputs_0 ? 7'h0 : _GEN_1500; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1502 = 10'h1de == io_inputs_0 ? 7'h0 : _GEN_1501; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1503 = 10'h1df == io_inputs_0 ? 7'h0 : _GEN_1502; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1504 = 10'h1e0 == io_inputs_0 ? 7'h0 : _GEN_1503; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1505 = 10'h1e1 == io_inputs_0 ? 7'h0 : _GEN_1504; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1506 = 10'h1e2 == io_inputs_0 ? 7'h0 : _GEN_1505; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1507 = 10'h1e3 == io_inputs_0 ? 7'h0 : _GEN_1506; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1508 = 10'h1e4 == io_inputs_0 ? 7'h0 : _GEN_1507; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1509 = 10'h1e5 == io_inputs_0 ? 7'h0 : _GEN_1508; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1510 = 10'h1e6 == io_inputs_0 ? 7'h0 : _GEN_1509; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1511 = 10'h1e7 == io_inputs_0 ? 7'h0 : _GEN_1510; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1512 = 10'h1e8 == io_inputs_0 ? 7'h0 : _GEN_1511; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1513 = 10'h1e9 == io_inputs_0 ? 7'h0 : _GEN_1512; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1514 = 10'h1ea == io_inputs_0 ? 7'h0 : _GEN_1513; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1515 = 10'h1eb == io_inputs_0 ? 7'h0 : _GEN_1514; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1516 = 10'h1ec == io_inputs_0 ? 7'h0 : _GEN_1515; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1517 = 10'h1ed == io_inputs_0 ? 7'h0 : _GEN_1516; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1518 = 10'h1ee == io_inputs_0 ? 7'h0 : _GEN_1517; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1519 = 10'h1ef == io_inputs_0 ? 7'h0 : _GEN_1518; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1520 = 10'h1f0 == io_inputs_0 ? 7'h0 : _GEN_1519; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1521 = 10'h1f1 == io_inputs_0 ? 7'h0 : _GEN_1520; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1522 = 10'h1f2 == io_inputs_0 ? 7'h0 : _GEN_1521; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1523 = 10'h1f3 == io_inputs_0 ? 7'h0 : _GEN_1522; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1524 = 10'h1f4 == io_inputs_0 ? 7'h0 : _GEN_1523; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1525 = 10'h1f5 == io_inputs_0 ? 7'h0 : _GEN_1524; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1526 = 10'h1f6 == io_inputs_0 ? 7'h0 : _GEN_1525; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1527 = 10'h1f7 == io_inputs_0 ? 7'h0 : _GEN_1526; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1528 = 10'h1f8 == io_inputs_0 ? 7'h0 : _GEN_1527; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1529 = 10'h1f9 == io_inputs_0 ? 7'h0 : _GEN_1528; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1530 = 10'h1fa == io_inputs_0 ? 7'h0 : _GEN_1529; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1531 = 10'h1fb == io_inputs_0 ? 7'h0 : _GEN_1530; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1532 = 10'h1fc == io_inputs_0 ? 7'h0 : _GEN_1531; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1533 = 10'h1fd == io_inputs_0 ? 7'h0 : _GEN_1532; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1534 = 10'h1fe == io_inputs_0 ? 7'h0 : _GEN_1533; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1535 = 10'h1ff == io_inputs_0 ? 7'h0 : _GEN_1534; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1536 = 10'h200 == io_inputs_0 ? 7'h0 : _GEN_1535; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1537 = 10'h201 == io_inputs_0 ? 7'h0 : _GEN_1536; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1538 = 10'h202 == io_inputs_0 ? 7'h0 : _GEN_1537; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1539 = 10'h203 == io_inputs_0 ? 7'h0 : _GEN_1538; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1540 = 10'h204 == io_inputs_0 ? 7'h0 : _GEN_1539; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1541 = 10'h205 == io_inputs_0 ? 7'h0 : _GEN_1540; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1542 = 10'h206 == io_inputs_0 ? 7'h0 : _GEN_1541; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1543 = 10'h207 == io_inputs_0 ? 7'h0 : _GEN_1542; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1544 = 10'h208 == io_inputs_0 ? 7'h0 : _GEN_1543; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1545 = 10'h209 == io_inputs_0 ? 7'h0 : _GEN_1544; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1546 = 10'h20a == io_inputs_0 ? 7'h0 : _GEN_1545; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1547 = 10'h20b == io_inputs_0 ? 7'h0 : _GEN_1546; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1548 = 10'h20c == io_inputs_0 ? 7'h0 : _GEN_1547; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1549 = 10'h20d == io_inputs_0 ? 7'h0 : _GEN_1548; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1550 = 10'h20e == io_inputs_0 ? 7'h0 : _GEN_1549; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1551 = 10'h20f == io_inputs_0 ? 7'h0 : _GEN_1550; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1552 = 10'h210 == io_inputs_0 ? 7'h0 : _GEN_1551; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1553 = 10'h211 == io_inputs_0 ? 7'h0 : _GEN_1552; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1554 = 10'h212 == io_inputs_0 ? 7'h0 : _GEN_1553; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1555 = 10'h213 == io_inputs_0 ? 7'h0 : _GEN_1554; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1556 = 10'h214 == io_inputs_0 ? 7'h0 : _GEN_1555; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1557 = 10'h215 == io_inputs_0 ? 7'h0 : _GEN_1556; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1558 = 10'h216 == io_inputs_0 ? 7'h0 : _GEN_1557; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1559 = 10'h217 == io_inputs_0 ? 7'h0 : _GEN_1558; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1560 = 10'h218 == io_inputs_0 ? 7'h0 : _GEN_1559; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1561 = 10'h219 == io_inputs_0 ? 7'h0 : _GEN_1560; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1562 = 10'h21a == io_inputs_0 ? 7'h0 : _GEN_1561; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1563 = 10'h21b == io_inputs_0 ? 7'h0 : _GEN_1562; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1564 = 10'h21c == io_inputs_0 ? 7'h0 : _GEN_1563; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1565 = 10'h21d == io_inputs_0 ? 7'h0 : _GEN_1564; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1566 = 10'h21e == io_inputs_0 ? 7'h0 : _GEN_1565; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1567 = 10'h21f == io_inputs_0 ? 7'h0 : _GEN_1566; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1568 = 10'h220 == io_inputs_0 ? 7'h0 : _GEN_1567; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1569 = 10'h221 == io_inputs_0 ? 7'h0 : _GEN_1568; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1570 = 10'h222 == io_inputs_0 ? 7'h0 : _GEN_1569; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1571 = 10'h223 == io_inputs_0 ? 7'h0 : _GEN_1570; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1572 = 10'h224 == io_inputs_0 ? 7'h0 : _GEN_1571; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1573 = 10'h225 == io_inputs_0 ? 7'h0 : _GEN_1572; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1574 = 10'h226 == io_inputs_0 ? 7'h0 : _GEN_1573; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1575 = 10'h227 == io_inputs_0 ? 7'h0 : _GEN_1574; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1576 = 10'h228 == io_inputs_0 ? 7'h0 : _GEN_1575; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1577 = 10'h229 == io_inputs_0 ? 7'h0 : _GEN_1576; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1578 = 10'h22a == io_inputs_0 ? 7'h0 : _GEN_1577; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1579 = 10'h22b == io_inputs_0 ? 7'h0 : _GEN_1578; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1580 = 10'h22c == io_inputs_0 ? 7'h0 : _GEN_1579; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1581 = 10'h22d == io_inputs_0 ? 7'h0 : _GEN_1580; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1582 = 10'h22e == io_inputs_0 ? 7'h0 : _GEN_1581; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1583 = 10'h22f == io_inputs_0 ? 7'h0 : _GEN_1582; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1584 = 10'h230 == io_inputs_0 ? 7'h0 : _GEN_1583; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1585 = 10'h231 == io_inputs_0 ? 7'h0 : _GEN_1584; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1586 = 10'h232 == io_inputs_0 ? 7'h0 : _GEN_1585; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1587 = 10'h233 == io_inputs_0 ? 7'h0 : _GEN_1586; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1588 = 10'h234 == io_inputs_0 ? 7'h0 : _GEN_1587; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1589 = 10'h235 == io_inputs_0 ? 7'h0 : _GEN_1588; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1590 = 10'h236 == io_inputs_0 ? 7'h0 : _GEN_1589; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1591 = 10'h237 == io_inputs_0 ? 7'h0 : _GEN_1590; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1592 = 10'h238 == io_inputs_0 ? 7'h0 : _GEN_1591; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1593 = 10'h239 == io_inputs_0 ? 7'h0 : _GEN_1592; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1594 = 10'h23a == io_inputs_0 ? 7'h0 : _GEN_1593; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1595 = 10'h23b == io_inputs_0 ? 7'h0 : _GEN_1594; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1596 = 10'h23c == io_inputs_0 ? 7'h0 : _GEN_1595; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1597 = 10'h23d == io_inputs_0 ? 7'h0 : _GEN_1596; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1598 = 10'h23e == io_inputs_0 ? 7'h0 : _GEN_1597; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1599 = 10'h23f == io_inputs_0 ? 7'h0 : _GEN_1598; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1600 = 10'h240 == io_inputs_0 ? 7'h0 : _GEN_1599; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1601 = 10'h241 == io_inputs_0 ? 7'h0 : _GEN_1600; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1602 = 10'h242 == io_inputs_0 ? 7'h0 : _GEN_1601; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1603 = 10'h243 == io_inputs_0 ? 7'h0 : _GEN_1602; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1604 = 10'h244 == io_inputs_0 ? 7'h0 : _GEN_1603; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1605 = 10'h245 == io_inputs_0 ? 7'h0 : _GEN_1604; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1606 = 10'h246 == io_inputs_0 ? 7'h0 : _GEN_1605; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1607 = 10'h247 == io_inputs_0 ? 7'h0 : _GEN_1606; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1608 = 10'h248 == io_inputs_0 ? 7'h0 : _GEN_1607; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1609 = 10'h249 == io_inputs_0 ? 7'h0 : _GEN_1608; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1610 = 10'h24a == io_inputs_0 ? 7'h0 : _GEN_1609; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1611 = 10'h24b == io_inputs_0 ? 7'h0 : _GEN_1610; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1612 = 10'h24c == io_inputs_0 ? 7'h0 : _GEN_1611; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1613 = 10'h24d == io_inputs_0 ? 7'h0 : _GEN_1612; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1614 = 10'h24e == io_inputs_0 ? 7'h0 : _GEN_1613; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1615 = 10'h24f == io_inputs_0 ? 7'h0 : _GEN_1614; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1616 = 10'h250 == io_inputs_0 ? 7'h0 : _GEN_1615; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1617 = 10'h251 == io_inputs_0 ? 7'h0 : _GEN_1616; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1618 = 10'h252 == io_inputs_0 ? 7'h0 : _GEN_1617; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1619 = 10'h253 == io_inputs_0 ? 7'h0 : _GEN_1618; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1620 = 10'h254 == io_inputs_0 ? 7'h0 : _GEN_1619; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1621 = 10'h255 == io_inputs_0 ? 7'h0 : _GEN_1620; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1622 = 10'h256 == io_inputs_0 ? 7'h0 : _GEN_1621; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1623 = 10'h257 == io_inputs_0 ? 7'h0 : _GEN_1622; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1624 = 10'h258 == io_inputs_0 ? 7'h0 : _GEN_1623; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1625 = 10'h259 == io_inputs_0 ? 7'h0 : _GEN_1624; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1626 = 10'h25a == io_inputs_0 ? 7'h0 : _GEN_1625; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1627 = 10'h25b == io_inputs_0 ? 7'h0 : _GEN_1626; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1628 = 10'h25c == io_inputs_0 ? 7'h0 : _GEN_1627; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1629 = 10'h25d == io_inputs_0 ? 7'h0 : _GEN_1628; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1630 = 10'h25e == io_inputs_0 ? 7'h0 : _GEN_1629; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1631 = 10'h25f == io_inputs_0 ? 7'h0 : _GEN_1630; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1632 = 10'h260 == io_inputs_0 ? 7'h0 : _GEN_1631; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1633 = 10'h261 == io_inputs_0 ? 7'h0 : _GEN_1632; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1634 = 10'h262 == io_inputs_0 ? 7'h0 : _GEN_1633; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1635 = 10'h263 == io_inputs_0 ? 7'h0 : _GEN_1634; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1636 = 10'h264 == io_inputs_0 ? 7'h0 : _GEN_1635; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1637 = 10'h265 == io_inputs_0 ? 7'h0 : _GEN_1636; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1638 = 10'h266 == io_inputs_0 ? 7'h0 : _GEN_1637; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1639 = 10'h267 == io_inputs_0 ? 7'h0 : _GEN_1638; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1640 = 10'h268 == io_inputs_0 ? 7'h0 : _GEN_1639; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1641 = 10'h269 == io_inputs_0 ? 7'h0 : _GEN_1640; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1642 = 10'h26a == io_inputs_0 ? 7'h0 : _GEN_1641; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1643 = 10'h26b == io_inputs_0 ? 7'h0 : _GEN_1642; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1644 = 10'h26c == io_inputs_0 ? 7'h0 : _GEN_1643; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1645 = 10'h26d == io_inputs_0 ? 7'h0 : _GEN_1644; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1646 = 10'h26e == io_inputs_0 ? 7'h0 : _GEN_1645; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1647 = 10'h26f == io_inputs_0 ? 7'h0 : _GEN_1646; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1648 = 10'h270 == io_inputs_0 ? 7'h0 : _GEN_1647; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1649 = 10'h271 == io_inputs_0 ? 7'h0 : _GEN_1648; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1650 = 10'h272 == io_inputs_0 ? 7'h0 : _GEN_1649; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1651 = 10'h273 == io_inputs_0 ? 7'h0 : _GEN_1650; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1652 = 10'h274 == io_inputs_0 ? 7'h0 : _GEN_1651; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1653 = 10'h275 == io_inputs_0 ? 7'h0 : _GEN_1652; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1654 = 10'h276 == io_inputs_0 ? 7'h0 : _GEN_1653; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1655 = 10'h277 == io_inputs_0 ? 7'h0 : _GEN_1654; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1656 = 10'h278 == io_inputs_0 ? 7'h0 : _GEN_1655; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1657 = 10'h279 == io_inputs_0 ? 7'h0 : _GEN_1656; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1658 = 10'h27a == io_inputs_0 ? 7'h0 : _GEN_1657; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1659 = 10'h27b == io_inputs_0 ? 7'h0 : _GEN_1658; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1660 = 10'h27c == io_inputs_0 ? 7'h0 : _GEN_1659; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1661 = 10'h27d == io_inputs_0 ? 7'h0 : _GEN_1660; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1662 = 10'h27e == io_inputs_0 ? 7'h0 : _GEN_1661; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1663 = 10'h27f == io_inputs_0 ? 7'h0 : _GEN_1662; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1664 = 10'h280 == io_inputs_0 ? 7'h0 : _GEN_1663; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1665 = 10'h281 == io_inputs_0 ? 7'h0 : _GEN_1664; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1666 = 10'h282 == io_inputs_0 ? 7'h0 : _GEN_1665; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1667 = 10'h283 == io_inputs_0 ? 7'h0 : _GEN_1666; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1668 = 10'h284 == io_inputs_0 ? 7'h0 : _GEN_1667; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1669 = 10'h285 == io_inputs_0 ? 7'h0 : _GEN_1668; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1670 = 10'h286 == io_inputs_0 ? 7'h0 : _GEN_1669; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1671 = 10'h287 == io_inputs_0 ? 7'h0 : _GEN_1670; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1672 = 10'h288 == io_inputs_0 ? 7'h0 : _GEN_1671; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1673 = 10'h289 == io_inputs_0 ? 7'h0 : _GEN_1672; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1674 = 10'h28a == io_inputs_0 ? 7'h0 : _GEN_1673; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1675 = 10'h28b == io_inputs_0 ? 7'h0 : _GEN_1674; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1676 = 10'h28c == io_inputs_0 ? 7'h0 : _GEN_1675; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1677 = 10'h28d == io_inputs_0 ? 7'h0 : _GEN_1676; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1678 = 10'h28e == io_inputs_0 ? 7'h0 : _GEN_1677; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1679 = 10'h28f == io_inputs_0 ? 7'h0 : _GEN_1678; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1680 = 10'h290 == io_inputs_0 ? 7'h0 : _GEN_1679; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1681 = 10'h291 == io_inputs_0 ? 7'h0 : _GEN_1680; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1682 = 10'h292 == io_inputs_0 ? 7'h0 : _GEN_1681; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1683 = 10'h293 == io_inputs_0 ? 7'h0 : _GEN_1682; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1684 = 10'h294 == io_inputs_0 ? 7'h0 : _GEN_1683; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1685 = 10'h295 == io_inputs_0 ? 7'h0 : _GEN_1684; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1686 = 10'h296 == io_inputs_0 ? 7'h0 : _GEN_1685; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1687 = 10'h297 == io_inputs_0 ? 7'h0 : _GEN_1686; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1688 = 10'h298 == io_inputs_0 ? 7'h0 : _GEN_1687; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1689 = 10'h299 == io_inputs_0 ? 7'h0 : _GEN_1688; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1690 = 10'h29a == io_inputs_0 ? 7'h0 : _GEN_1689; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1691 = 10'h29b == io_inputs_0 ? 7'h0 : _GEN_1690; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1692 = 10'h29c == io_inputs_0 ? 7'h0 : _GEN_1691; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1693 = 10'h29d == io_inputs_0 ? 7'h0 : _GEN_1692; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1694 = 10'h29e == io_inputs_0 ? 7'h0 : _GEN_1693; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1695 = 10'h29f == io_inputs_0 ? 7'h0 : _GEN_1694; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1696 = 10'h2a0 == io_inputs_0 ? 7'h0 : _GEN_1695; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1697 = 10'h2a1 == io_inputs_0 ? 7'h0 : _GEN_1696; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1698 = 10'h2a2 == io_inputs_0 ? 7'h0 : _GEN_1697; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1699 = 10'h2a3 == io_inputs_0 ? 7'h0 : _GEN_1698; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1700 = 10'h2a4 == io_inputs_0 ? 7'h0 : _GEN_1699; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1701 = 10'h2a5 == io_inputs_0 ? 7'h0 : _GEN_1700; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1702 = 10'h2a6 == io_inputs_0 ? 7'h0 : _GEN_1701; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1703 = 10'h2a7 == io_inputs_0 ? 7'h0 : _GEN_1702; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1704 = 10'h2a8 == io_inputs_0 ? 7'h0 : _GEN_1703; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1705 = 10'h2a9 == io_inputs_0 ? 7'h0 : _GEN_1704; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1706 = 10'h2aa == io_inputs_0 ? 7'h0 : _GEN_1705; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1707 = 10'h2ab == io_inputs_0 ? 7'h0 : _GEN_1706; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1708 = 10'h2ac == io_inputs_0 ? 7'h0 : _GEN_1707; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1709 = 10'h2ad == io_inputs_0 ? 7'h0 : _GEN_1708; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1710 = 10'h2ae == io_inputs_0 ? 7'h0 : _GEN_1709; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1711 = 10'h2af == io_inputs_0 ? 7'h0 : _GEN_1710; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1712 = 10'h2b0 == io_inputs_0 ? 7'h0 : _GEN_1711; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1713 = 10'h2b1 == io_inputs_0 ? 7'h0 : _GEN_1712; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1714 = 10'h2b2 == io_inputs_0 ? 7'h0 : _GEN_1713; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1715 = 10'h2b3 == io_inputs_0 ? 7'h0 : _GEN_1714; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1716 = 10'h2b4 == io_inputs_0 ? 7'h0 : _GEN_1715; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1717 = 10'h2b5 == io_inputs_0 ? 7'h0 : _GEN_1716; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1718 = 10'h2b6 == io_inputs_0 ? 7'h0 : _GEN_1717; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1719 = 10'h2b7 == io_inputs_0 ? 7'h0 : _GEN_1718; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1720 = 10'h2b8 == io_inputs_0 ? 7'h0 : _GEN_1719; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1721 = 10'h2b9 == io_inputs_0 ? 7'h0 : _GEN_1720; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1722 = 10'h2ba == io_inputs_0 ? 7'h0 : _GEN_1721; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1723 = 10'h2bb == io_inputs_0 ? 7'h0 : _GEN_1722; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1724 = 10'h2bc == io_inputs_0 ? 7'h0 : _GEN_1723; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1725 = 10'h2bd == io_inputs_0 ? 7'h0 : _GEN_1724; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1726 = 10'h2be == io_inputs_0 ? 7'h0 : _GEN_1725; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1727 = 10'h2bf == io_inputs_0 ? 7'h0 : _GEN_1726; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1728 = 10'h2c0 == io_inputs_0 ? 7'h0 : _GEN_1727; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1729 = 10'h2c1 == io_inputs_0 ? 7'h0 : _GEN_1728; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1730 = 10'h2c2 == io_inputs_0 ? 7'h0 : _GEN_1729; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1731 = 10'h2c3 == io_inputs_0 ? 7'h0 : _GEN_1730; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1732 = 10'h2c4 == io_inputs_0 ? 7'h0 : _GEN_1731; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1733 = 10'h2c5 == io_inputs_0 ? 7'h0 : _GEN_1732; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1734 = 10'h2c6 == io_inputs_0 ? 7'h0 : _GEN_1733; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1735 = 10'h2c7 == io_inputs_0 ? 7'h0 : _GEN_1734; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1736 = 10'h2c8 == io_inputs_0 ? 7'h0 : _GEN_1735; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1737 = 10'h2c9 == io_inputs_0 ? 7'h0 : _GEN_1736; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1738 = 10'h2ca == io_inputs_0 ? 7'h0 : _GEN_1737; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1739 = 10'h2cb == io_inputs_0 ? 7'h0 : _GEN_1738; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1740 = 10'h2cc == io_inputs_0 ? 7'h0 : _GEN_1739; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1741 = 10'h2cd == io_inputs_0 ? 7'h0 : _GEN_1740; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1742 = 10'h2ce == io_inputs_0 ? 7'h0 : _GEN_1741; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1743 = 10'h2cf == io_inputs_0 ? 7'h0 : _GEN_1742; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1744 = 10'h2d0 == io_inputs_0 ? 7'h0 : _GEN_1743; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1745 = 10'h2d1 == io_inputs_0 ? 7'h0 : _GEN_1744; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1746 = 10'h2d2 == io_inputs_0 ? 7'h0 : _GEN_1745; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1747 = 10'h2d3 == io_inputs_0 ? 7'h0 : _GEN_1746; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1748 = 10'h2d4 == io_inputs_0 ? 7'h0 : _GEN_1747; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1749 = 10'h2d5 == io_inputs_0 ? 7'h0 : _GEN_1748; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1750 = 10'h2d6 == io_inputs_0 ? 7'h0 : _GEN_1749; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1751 = 10'h2d7 == io_inputs_0 ? 7'h0 : _GEN_1750; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1752 = 10'h2d8 == io_inputs_0 ? 7'h0 : _GEN_1751; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1753 = 10'h2d9 == io_inputs_0 ? 7'h0 : _GEN_1752; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1754 = 10'h2da == io_inputs_0 ? 7'h0 : _GEN_1753; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1755 = 10'h2db == io_inputs_0 ? 7'h0 : _GEN_1754; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1756 = 10'h2dc == io_inputs_0 ? 7'h0 : _GEN_1755; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1757 = 10'h2dd == io_inputs_0 ? 7'h0 : _GEN_1756; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1758 = 10'h2de == io_inputs_0 ? 7'h0 : _GEN_1757; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1759 = 10'h2df == io_inputs_0 ? 7'h0 : _GEN_1758; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1760 = 10'h2e0 == io_inputs_0 ? 7'h0 : _GEN_1759; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1761 = 10'h2e1 == io_inputs_0 ? 7'h0 : _GEN_1760; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1762 = 10'h2e2 == io_inputs_0 ? 7'h0 : _GEN_1761; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1763 = 10'h2e3 == io_inputs_0 ? 7'h0 : _GEN_1762; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1764 = 10'h2e4 == io_inputs_0 ? 7'h0 : _GEN_1763; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1765 = 10'h2e5 == io_inputs_0 ? 7'h0 : _GEN_1764; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1766 = 10'h2e6 == io_inputs_0 ? 7'h0 : _GEN_1765; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1767 = 10'h2e7 == io_inputs_0 ? 7'h0 : _GEN_1766; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1768 = 10'h2e8 == io_inputs_0 ? 7'h0 : _GEN_1767; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1769 = 10'h2e9 == io_inputs_0 ? 7'h0 : _GEN_1768; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1770 = 10'h2ea == io_inputs_0 ? 7'h0 : _GEN_1769; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1771 = 10'h2eb == io_inputs_0 ? 7'h0 : _GEN_1770; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1772 = 10'h2ec == io_inputs_0 ? 7'h0 : _GEN_1771; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1773 = 10'h2ed == io_inputs_0 ? 7'h0 : _GEN_1772; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1774 = 10'h2ee == io_inputs_0 ? 7'h0 : _GEN_1773; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1775 = 10'h2ef == io_inputs_0 ? 7'h0 : _GEN_1774; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1776 = 10'h2f0 == io_inputs_0 ? 7'h0 : _GEN_1775; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1777 = 10'h2f1 == io_inputs_0 ? 7'h0 : _GEN_1776; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1778 = 10'h2f2 == io_inputs_0 ? 7'h0 : _GEN_1777; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1779 = 10'h2f3 == io_inputs_0 ? 7'h0 : _GEN_1778; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1780 = 10'h2f4 == io_inputs_0 ? 7'h0 : _GEN_1779; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1781 = 10'h2f5 == io_inputs_0 ? 7'h0 : _GEN_1780; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1782 = 10'h2f6 == io_inputs_0 ? 7'h0 : _GEN_1781; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1783 = 10'h2f7 == io_inputs_0 ? 7'h0 : _GEN_1782; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1784 = 10'h2f8 == io_inputs_0 ? 7'h0 : _GEN_1783; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1785 = 10'h2f9 == io_inputs_0 ? 7'h0 : _GEN_1784; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1786 = 10'h2fa == io_inputs_0 ? 7'h0 : _GEN_1785; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1787 = 10'h2fb == io_inputs_0 ? 7'h0 : _GEN_1786; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1788 = 10'h2fc == io_inputs_0 ? 7'h0 : _GEN_1787; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1789 = 10'h2fd == io_inputs_0 ? 7'h0 : _GEN_1788; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1790 = 10'h2fe == io_inputs_0 ? 7'h0 : _GEN_1789; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1791 = 10'h2ff == io_inputs_0 ? 7'h0 : _GEN_1790; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1792 = 10'h300 == io_inputs_0 ? 7'h0 : _GEN_1791; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1793 = 10'h301 == io_inputs_0 ? 7'h0 : _GEN_1792; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1794 = 10'h302 == io_inputs_0 ? 7'h0 : _GEN_1793; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1795 = 10'h303 == io_inputs_0 ? 7'h0 : _GEN_1794; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1796 = 10'h304 == io_inputs_0 ? 7'h0 : _GEN_1795; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1797 = 10'h305 == io_inputs_0 ? 7'h0 : _GEN_1796; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1798 = 10'h306 == io_inputs_0 ? 7'h0 : _GEN_1797; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1799 = 10'h307 == io_inputs_0 ? 7'h0 : _GEN_1798; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1800 = 10'h308 == io_inputs_0 ? 7'h0 : _GEN_1799; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1801 = 10'h309 == io_inputs_0 ? 7'h0 : _GEN_1800; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1802 = 10'h30a == io_inputs_0 ? 7'h0 : _GEN_1801; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1803 = 10'h30b == io_inputs_0 ? 7'h0 : _GEN_1802; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1804 = 10'h30c == io_inputs_0 ? 7'h0 : _GEN_1803; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1805 = 10'h30d == io_inputs_0 ? 7'h0 : _GEN_1804; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1806 = 10'h30e == io_inputs_0 ? 7'h0 : _GEN_1805; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1807 = 10'h30f == io_inputs_0 ? 7'h0 : _GEN_1806; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1808 = 10'h310 == io_inputs_0 ? 7'h0 : _GEN_1807; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1809 = 10'h311 == io_inputs_0 ? 7'h0 : _GEN_1808; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1810 = 10'h312 == io_inputs_0 ? 7'h0 : _GEN_1809; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1811 = 10'h313 == io_inputs_0 ? 7'h0 : _GEN_1810; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1812 = 10'h314 == io_inputs_0 ? 7'h0 : _GEN_1811; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1813 = 10'h315 == io_inputs_0 ? 7'h0 : _GEN_1812; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1814 = 10'h316 == io_inputs_0 ? 7'h0 : _GEN_1813; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1815 = 10'h317 == io_inputs_0 ? 7'h0 : _GEN_1814; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1816 = 10'h318 == io_inputs_0 ? 7'h0 : _GEN_1815; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1817 = 10'h319 == io_inputs_0 ? 7'h0 : _GEN_1816; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1818 = 10'h31a == io_inputs_0 ? 7'h0 : _GEN_1817; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1819 = 10'h31b == io_inputs_0 ? 7'h0 : _GEN_1818; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1820 = 10'h31c == io_inputs_0 ? 7'h0 : _GEN_1819; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1821 = 10'h31d == io_inputs_0 ? 7'h0 : _GEN_1820; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1822 = 10'h31e == io_inputs_0 ? 7'h0 : _GEN_1821; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1823 = 10'h31f == io_inputs_0 ? 7'h0 : _GEN_1822; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1824 = 10'h320 == io_inputs_0 ? 7'h0 : _GEN_1823; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1825 = 10'h321 == io_inputs_0 ? 7'h0 : _GEN_1824; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1826 = 10'h322 == io_inputs_0 ? 7'h0 : _GEN_1825; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1827 = 10'h323 == io_inputs_0 ? 7'h0 : _GEN_1826; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1828 = 10'h324 == io_inputs_0 ? 7'h0 : _GEN_1827; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1829 = 10'h325 == io_inputs_0 ? 7'h0 : _GEN_1828; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1830 = 10'h326 == io_inputs_0 ? 7'h0 : _GEN_1829; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1831 = 10'h327 == io_inputs_0 ? 7'h0 : _GEN_1830; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1832 = 10'h328 == io_inputs_0 ? 7'h0 : _GEN_1831; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1833 = 10'h329 == io_inputs_0 ? 7'h0 : _GEN_1832; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1834 = 10'h32a == io_inputs_0 ? 7'h0 : _GEN_1833; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1835 = 10'h32b == io_inputs_0 ? 7'h0 : _GEN_1834; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1836 = 10'h32c == io_inputs_0 ? 7'h0 : _GEN_1835; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1837 = 10'h32d == io_inputs_0 ? 7'h0 : _GEN_1836; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1838 = 10'h32e == io_inputs_0 ? 7'h0 : _GEN_1837; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1839 = 10'h32f == io_inputs_0 ? 7'h0 : _GEN_1838; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1840 = 10'h330 == io_inputs_0 ? 7'h0 : _GEN_1839; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1841 = 10'h331 == io_inputs_0 ? 7'h0 : _GEN_1840; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1842 = 10'h332 == io_inputs_0 ? 7'h0 : _GEN_1841; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1843 = 10'h333 == io_inputs_0 ? 7'h0 : _GEN_1842; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1844 = 10'h334 == io_inputs_0 ? 7'h0 : _GEN_1843; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1845 = 10'h335 == io_inputs_0 ? 7'h0 : _GEN_1844; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1846 = 10'h336 == io_inputs_0 ? 7'h0 : _GEN_1845; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1847 = 10'h337 == io_inputs_0 ? 7'h0 : _GEN_1846; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1848 = 10'h338 == io_inputs_0 ? 7'h0 : _GEN_1847; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1849 = 10'h339 == io_inputs_0 ? 7'h0 : _GEN_1848; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1850 = 10'h33a == io_inputs_0 ? 7'h0 : _GEN_1849; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1851 = 10'h33b == io_inputs_0 ? 7'h0 : _GEN_1850; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1852 = 10'h33c == io_inputs_0 ? 7'h0 : _GEN_1851; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1853 = 10'h33d == io_inputs_0 ? 7'h0 : _GEN_1852; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1854 = 10'h33e == io_inputs_0 ? 7'h0 : _GEN_1853; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1855 = 10'h33f == io_inputs_0 ? 7'h0 : _GEN_1854; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1856 = 10'h340 == io_inputs_0 ? 7'h0 : _GEN_1855; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1857 = 10'h341 == io_inputs_0 ? 7'h0 : _GEN_1856; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1858 = 10'h342 == io_inputs_0 ? 7'h0 : _GEN_1857; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1859 = 10'h343 == io_inputs_0 ? 7'h0 : _GEN_1858; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1860 = 10'h344 == io_inputs_0 ? 7'h0 : _GEN_1859; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1861 = 10'h345 == io_inputs_0 ? 7'h0 : _GEN_1860; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1862 = 10'h346 == io_inputs_0 ? 7'h0 : _GEN_1861; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1863 = 10'h347 == io_inputs_0 ? 7'h0 : _GEN_1862; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1864 = 10'h348 == io_inputs_0 ? 7'h0 : _GEN_1863; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1865 = 10'h349 == io_inputs_0 ? 7'h0 : _GEN_1864; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1866 = 10'h34a == io_inputs_0 ? 7'h0 : _GEN_1865; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1867 = 10'h34b == io_inputs_0 ? 7'h0 : _GEN_1866; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1868 = 10'h34c == io_inputs_0 ? 7'h0 : _GEN_1867; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1869 = 10'h34d == io_inputs_0 ? 7'h0 : _GEN_1868; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1870 = 10'h34e == io_inputs_0 ? 7'h0 : _GEN_1869; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1871 = 10'h34f == io_inputs_0 ? 7'h0 : _GEN_1870; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1872 = 10'h350 == io_inputs_0 ? 7'h0 : _GEN_1871; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1873 = 10'h351 == io_inputs_0 ? 7'h0 : _GEN_1872; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1874 = 10'h352 == io_inputs_0 ? 7'h0 : _GEN_1873; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1875 = 10'h353 == io_inputs_0 ? 7'h0 : _GEN_1874; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1876 = 10'h354 == io_inputs_0 ? 7'h0 : _GEN_1875; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1877 = 10'h355 == io_inputs_0 ? 7'h0 : _GEN_1876; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1878 = 10'h356 == io_inputs_0 ? 7'h0 : _GEN_1877; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1879 = 10'h357 == io_inputs_0 ? 7'h0 : _GEN_1878; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1880 = 10'h358 == io_inputs_0 ? 7'h0 : _GEN_1879; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1881 = 10'h359 == io_inputs_0 ? 7'h0 : _GEN_1880; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1882 = 10'h35a == io_inputs_0 ? 7'h0 : _GEN_1881; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1883 = 10'h35b == io_inputs_0 ? 7'h0 : _GEN_1882; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1884 = 10'h35c == io_inputs_0 ? 7'h0 : _GEN_1883; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1885 = 10'h35d == io_inputs_0 ? 7'h0 : _GEN_1884; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1886 = 10'h35e == io_inputs_0 ? 7'h0 : _GEN_1885; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1887 = 10'h35f == io_inputs_0 ? 7'h0 : _GEN_1886; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1888 = 10'h360 == io_inputs_0 ? 7'h0 : _GEN_1887; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1889 = 10'h361 == io_inputs_0 ? 7'h0 : _GEN_1888; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1890 = 10'h362 == io_inputs_0 ? 7'h0 : _GEN_1889; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1891 = 10'h363 == io_inputs_0 ? 7'h0 : _GEN_1890; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1892 = 10'h364 == io_inputs_0 ? 7'h0 : _GEN_1891; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1893 = 10'h365 == io_inputs_0 ? 7'h0 : _GEN_1892; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1894 = 10'h366 == io_inputs_0 ? 7'h0 : _GEN_1893; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1895 = 10'h367 == io_inputs_0 ? 7'h0 : _GEN_1894; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1896 = 10'h368 == io_inputs_0 ? 7'h0 : _GEN_1895; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1897 = 10'h369 == io_inputs_0 ? 7'h0 : _GEN_1896; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1898 = 10'h36a == io_inputs_0 ? 7'h0 : _GEN_1897; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1899 = 10'h36b == io_inputs_0 ? 7'h0 : _GEN_1898; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1900 = 10'h36c == io_inputs_0 ? 7'h0 : _GEN_1899; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1901 = 10'h36d == io_inputs_0 ? 7'h0 : _GEN_1900; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1902 = 10'h36e == io_inputs_0 ? 7'h0 : _GEN_1901; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1903 = 10'h36f == io_inputs_0 ? 7'h0 : _GEN_1902; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1904 = 10'h370 == io_inputs_0 ? 7'h0 : _GEN_1903; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1905 = 10'h371 == io_inputs_0 ? 7'h0 : _GEN_1904; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1906 = 10'h372 == io_inputs_0 ? 7'h0 : _GEN_1905; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1907 = 10'h373 == io_inputs_0 ? 7'h0 : _GEN_1906; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1908 = 10'h374 == io_inputs_0 ? 7'h0 : _GEN_1907; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1909 = 10'h375 == io_inputs_0 ? 7'h0 : _GEN_1908; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1910 = 10'h376 == io_inputs_0 ? 7'h0 : _GEN_1909; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1911 = 10'h377 == io_inputs_0 ? 7'h0 : _GEN_1910; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1912 = 10'h378 == io_inputs_0 ? 7'h0 : _GEN_1911; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1913 = 10'h379 == io_inputs_0 ? 7'h0 : _GEN_1912; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1914 = 10'h37a == io_inputs_0 ? 7'h0 : _GEN_1913; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1915 = 10'h37b == io_inputs_0 ? 7'h0 : _GEN_1914; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1916 = 10'h37c == io_inputs_0 ? 7'h0 : _GEN_1915; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1917 = 10'h37d == io_inputs_0 ? 7'h0 : _GEN_1916; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1918 = 10'h37e == io_inputs_0 ? 7'h0 : _GEN_1917; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1919 = 10'h37f == io_inputs_0 ? 7'h0 : _GEN_1918; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1920 = 10'h380 == io_inputs_0 ? 7'h0 : _GEN_1919; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1921 = 10'h381 == io_inputs_0 ? 7'h0 : _GEN_1920; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1922 = 10'h382 == io_inputs_0 ? 7'h0 : _GEN_1921; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1923 = 10'h383 == io_inputs_0 ? 7'h0 : _GEN_1922; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1924 = 10'h384 == io_inputs_0 ? 7'h0 : _GEN_1923; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1925 = 10'h385 == io_inputs_0 ? 7'h0 : _GEN_1924; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1926 = 10'h386 == io_inputs_0 ? 7'h0 : _GEN_1925; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1927 = 10'h387 == io_inputs_0 ? 7'h0 : _GEN_1926; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1928 = 10'h388 == io_inputs_0 ? 7'h0 : _GEN_1927; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1929 = 10'h389 == io_inputs_0 ? 7'h0 : _GEN_1928; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1930 = 10'h38a == io_inputs_0 ? 7'h0 : _GEN_1929; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1931 = 10'h38b == io_inputs_0 ? 7'h0 : _GEN_1930; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1932 = 10'h38c == io_inputs_0 ? 7'h0 : _GEN_1931; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1933 = 10'h38d == io_inputs_0 ? 7'h0 : _GEN_1932; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1934 = 10'h38e == io_inputs_0 ? 7'h0 : _GEN_1933; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1935 = 10'h38f == io_inputs_0 ? 7'h0 : _GEN_1934; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1936 = 10'h390 == io_inputs_0 ? 7'h0 : _GEN_1935; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1937 = 10'h391 == io_inputs_0 ? 7'h0 : _GEN_1936; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1938 = 10'h392 == io_inputs_0 ? 7'h0 : _GEN_1937; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1939 = 10'h393 == io_inputs_0 ? 7'h0 : _GEN_1938; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1940 = 10'h394 == io_inputs_0 ? 7'h0 : _GEN_1939; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1941 = 10'h395 == io_inputs_0 ? 7'h0 : _GEN_1940; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1942 = 10'h396 == io_inputs_0 ? 7'h0 : _GEN_1941; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1943 = 10'h397 == io_inputs_0 ? 7'h0 : _GEN_1942; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1944 = 10'h398 == io_inputs_0 ? 7'h0 : _GEN_1943; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1945 = 10'h399 == io_inputs_0 ? 7'h0 : _GEN_1944; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1946 = 10'h39a == io_inputs_0 ? 7'h0 : _GEN_1945; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1947 = 10'h39b == io_inputs_0 ? 7'h0 : _GEN_1946; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1948 = 10'h39c == io_inputs_0 ? 7'h0 : _GEN_1947; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1949 = 10'h39d == io_inputs_0 ? 7'h0 : _GEN_1948; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1950 = 10'h39e == io_inputs_0 ? 7'h0 : _GEN_1949; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1951 = 10'h39f == io_inputs_0 ? 7'h0 : _GEN_1950; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1952 = 10'h3a0 == io_inputs_0 ? 7'h0 : _GEN_1951; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1953 = 10'h3a1 == io_inputs_0 ? 7'h0 : _GEN_1952; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1954 = 10'h3a2 == io_inputs_0 ? 7'h0 : _GEN_1953; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1955 = 10'h3a3 == io_inputs_0 ? 7'h0 : _GEN_1954; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1956 = 10'h3a4 == io_inputs_0 ? 7'h0 : _GEN_1955; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1957 = 10'h3a5 == io_inputs_0 ? 7'h0 : _GEN_1956; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1958 = 10'h3a6 == io_inputs_0 ? 7'h0 : _GEN_1957; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1959 = 10'h3a7 == io_inputs_0 ? 7'h0 : _GEN_1958; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1960 = 10'h3a8 == io_inputs_0 ? 7'h0 : _GEN_1959; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1961 = 10'h3a9 == io_inputs_0 ? 7'h0 : _GEN_1960; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1962 = 10'h3aa == io_inputs_0 ? 7'h0 : _GEN_1961; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1963 = 10'h3ab == io_inputs_0 ? 7'h0 : _GEN_1962; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1964 = 10'h3ac == io_inputs_0 ? 7'h0 : _GEN_1963; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1965 = 10'h3ad == io_inputs_0 ? 7'h0 : _GEN_1964; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1966 = 10'h3ae == io_inputs_0 ? 7'h0 : _GEN_1965; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1967 = 10'h3af == io_inputs_0 ? 7'h0 : _GEN_1966; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1968 = 10'h3b0 == io_inputs_0 ? 7'h0 : _GEN_1967; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1969 = 10'h3b1 == io_inputs_0 ? 7'h0 : _GEN_1968; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1970 = 10'h3b2 == io_inputs_0 ? 7'h0 : _GEN_1969; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1971 = 10'h3b3 == io_inputs_0 ? 7'h0 : _GEN_1970; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1972 = 10'h3b4 == io_inputs_0 ? 7'h0 : _GEN_1971; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1973 = 10'h3b5 == io_inputs_0 ? 7'h0 : _GEN_1972; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1974 = 10'h3b6 == io_inputs_0 ? 7'h0 : _GEN_1973; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1975 = 10'h3b7 == io_inputs_0 ? 7'h0 : _GEN_1974; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1976 = 10'h3b8 == io_inputs_0 ? 7'h0 : _GEN_1975; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1977 = 10'h3b9 == io_inputs_0 ? 7'h0 : _GEN_1976; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1978 = 10'h3ba == io_inputs_0 ? 7'h0 : _GEN_1977; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1979 = 10'h3bb == io_inputs_0 ? 7'h0 : _GEN_1978; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1980 = 10'h3bc == io_inputs_0 ? 7'h0 : _GEN_1979; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1981 = 10'h3bd == io_inputs_0 ? 7'h0 : _GEN_1980; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1982 = 10'h3be == io_inputs_0 ? 7'h0 : _GEN_1981; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1983 = 10'h3bf == io_inputs_0 ? 7'h0 : _GEN_1982; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1984 = 10'h3c0 == io_inputs_0 ? 7'h0 : _GEN_1983; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1985 = 10'h3c1 == io_inputs_0 ? 7'h0 : _GEN_1984; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1986 = 10'h3c2 == io_inputs_0 ? 7'h0 : _GEN_1985; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1987 = 10'h3c3 == io_inputs_0 ? 7'h0 : _GEN_1986; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1988 = 10'h3c4 == io_inputs_0 ? 7'h0 : _GEN_1987; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1989 = 10'h3c5 == io_inputs_0 ? 7'h0 : _GEN_1988; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1990 = 10'h3c6 == io_inputs_0 ? 7'h0 : _GEN_1989; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1991 = 10'h3c7 == io_inputs_0 ? 7'h0 : _GEN_1990; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1992 = 10'h3c8 == io_inputs_0 ? 7'h0 : _GEN_1991; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1993 = 10'h3c9 == io_inputs_0 ? 7'h0 : _GEN_1992; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1994 = 10'h3ca == io_inputs_0 ? 7'h0 : _GEN_1993; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1995 = 10'h3cb == io_inputs_0 ? 7'h0 : _GEN_1994; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1996 = 10'h3cc == io_inputs_0 ? 7'h0 : _GEN_1995; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1997 = 10'h3cd == io_inputs_0 ? 7'h0 : _GEN_1996; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1998 = 10'h3ce == io_inputs_0 ? 7'h0 : _GEN_1997; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_1999 = 10'h3cf == io_inputs_0 ? 7'h0 : _GEN_1998; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2000 = 10'h3d0 == io_inputs_0 ? 7'h0 : _GEN_1999; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2001 = 10'h3d1 == io_inputs_0 ? 7'h0 : _GEN_2000; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2002 = 10'h3d2 == io_inputs_0 ? 7'h0 : _GEN_2001; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2003 = 10'h3d3 == io_inputs_0 ? 7'h0 : _GEN_2002; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2004 = 10'h3d4 == io_inputs_0 ? 7'h0 : _GEN_2003; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2005 = 10'h3d5 == io_inputs_0 ? 7'h0 : _GEN_2004; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2006 = 10'h3d6 == io_inputs_0 ? 7'h0 : _GEN_2005; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2007 = 10'h3d7 == io_inputs_0 ? 7'h0 : _GEN_2006; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2008 = 10'h3d8 == io_inputs_0 ? 7'h0 : _GEN_2007; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2009 = 10'h3d9 == io_inputs_0 ? 7'h0 : _GEN_2008; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2010 = 10'h3da == io_inputs_0 ? 7'h0 : _GEN_2009; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2011 = 10'h3db == io_inputs_0 ? 7'h0 : _GEN_2010; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2012 = 10'h3dc == io_inputs_0 ? 7'h0 : _GEN_2011; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2013 = 10'h3dd == io_inputs_0 ? 7'h0 : _GEN_2012; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2014 = 10'h3de == io_inputs_0 ? 7'h0 : _GEN_2013; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2015 = 10'h3df == io_inputs_0 ? 7'h0 : _GEN_2014; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2016 = 10'h3e0 == io_inputs_0 ? 7'h0 : _GEN_2015; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2017 = 10'h3e1 == io_inputs_0 ? 7'h0 : _GEN_2016; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2018 = 10'h3e2 == io_inputs_0 ? 7'h0 : _GEN_2017; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2019 = 10'h3e3 == io_inputs_0 ? 7'h0 : _GEN_2018; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2020 = 10'h3e4 == io_inputs_0 ? 7'h0 : _GEN_2019; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2021 = 10'h3e5 == io_inputs_0 ? 7'h0 : _GEN_2020; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2022 = 10'h3e6 == io_inputs_0 ? 7'h0 : _GEN_2021; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2023 = 10'h3e7 == io_inputs_0 ? 7'h0 : _GEN_2022; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2024 = 10'h3e8 == io_inputs_0 ? 7'h0 : _GEN_2023; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2025 = 10'h3e9 == io_inputs_0 ? 7'h0 : _GEN_2024; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2026 = 10'h3ea == io_inputs_0 ? 7'h0 : _GEN_2025; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2027 = 10'h3eb == io_inputs_0 ? 7'h0 : _GEN_2026; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2028 = 10'h3ec == io_inputs_0 ? 7'h0 : _GEN_2027; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2029 = 10'h3ed == io_inputs_0 ? 7'h0 : _GEN_2028; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2030 = 10'h3ee == io_inputs_0 ? 7'h0 : _GEN_2029; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2031 = 10'h3ef == io_inputs_0 ? 7'h0 : _GEN_2030; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2032 = 10'h3f0 == io_inputs_0 ? 7'h0 : _GEN_2031; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2033 = 10'h3f1 == io_inputs_0 ? 7'h0 : _GEN_2032; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2034 = 10'h3f2 == io_inputs_0 ? 7'h0 : _GEN_2033; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2035 = 10'h3f3 == io_inputs_0 ? 7'h0 : _GEN_2034; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2036 = 10'h3f4 == io_inputs_0 ? 7'h0 : _GEN_2035; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2037 = 10'h3f5 == io_inputs_0 ? 7'h0 : _GEN_2036; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2038 = 10'h3f6 == io_inputs_0 ? 7'h0 : _GEN_2037; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2039 = 10'h3f7 == io_inputs_0 ? 7'h0 : _GEN_2038; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2040 = 10'h3f8 == io_inputs_0 ? 7'h0 : _GEN_2039; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2041 = 10'h3f9 == io_inputs_0 ? 7'h0 : _GEN_2040; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2042 = 10'h3fa == io_inputs_0 ? 7'h0 : _GEN_2041; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2043 = 10'h3fb == io_inputs_0 ? 7'h0 : _GEN_2042; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2044 = 10'h3fc == io_inputs_0 ? 7'h0 : _GEN_2043; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2249 = 10'hc9 == io_inputs_0 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2250 = 10'hca == io_inputs_0 ? 7'h2 : _GEN_2249; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2251 = 10'hcb == io_inputs_0 ? 7'h3 : _GEN_2250; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2252 = 10'hcc == io_inputs_0 ? 7'h4 : _GEN_2251; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2253 = 10'hcd == io_inputs_0 ? 7'h5 : _GEN_2252; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2254 = 10'hce == io_inputs_0 ? 7'h6 : _GEN_2253; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2255 = 10'hcf == io_inputs_0 ? 7'h7 : _GEN_2254; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2256 = 10'hd0 == io_inputs_0 ? 7'h8 : _GEN_2255; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2257 = 10'hd1 == io_inputs_0 ? 7'h9 : _GEN_2256; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2258 = 10'hd2 == io_inputs_0 ? 7'ha : _GEN_2257; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2259 = 10'hd3 == io_inputs_0 ? 7'hb : _GEN_2258; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2260 = 10'hd4 == io_inputs_0 ? 7'hc : _GEN_2259; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2261 = 10'hd5 == io_inputs_0 ? 7'hd : _GEN_2260; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2262 = 10'hd6 == io_inputs_0 ? 7'he : _GEN_2261; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2263 = 10'hd7 == io_inputs_0 ? 7'hf : _GEN_2262; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2264 = 10'hd8 == io_inputs_0 ? 7'h10 : _GEN_2263; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2265 = 10'hd9 == io_inputs_0 ? 7'h11 : _GEN_2264; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2266 = 10'hda == io_inputs_0 ? 7'h12 : _GEN_2265; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2267 = 10'hdb == io_inputs_0 ? 7'h13 : _GEN_2266; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2268 = 10'hdc == io_inputs_0 ? 7'h14 : _GEN_2267; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2269 = 10'hdd == io_inputs_0 ? 7'h15 : _GEN_2268; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2270 = 10'hde == io_inputs_0 ? 7'h16 : _GEN_2269; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2271 = 10'hdf == io_inputs_0 ? 7'h17 : _GEN_2270; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2272 = 10'he0 == io_inputs_0 ? 7'h18 : _GEN_2271; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2273 = 10'he1 == io_inputs_0 ? 7'h19 : _GEN_2272; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2274 = 10'he2 == io_inputs_0 ? 7'h1a : _GEN_2273; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2275 = 10'he3 == io_inputs_0 ? 7'h1b : _GEN_2274; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2276 = 10'he4 == io_inputs_0 ? 7'h1c : _GEN_2275; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2277 = 10'he5 == io_inputs_0 ? 7'h1d : _GEN_2276; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2278 = 10'he6 == io_inputs_0 ? 7'h1e : _GEN_2277; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2279 = 10'he7 == io_inputs_0 ? 7'h1f : _GEN_2278; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2280 = 10'he8 == io_inputs_0 ? 7'h20 : _GEN_2279; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2281 = 10'he9 == io_inputs_0 ? 7'h21 : _GEN_2280; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2282 = 10'hea == io_inputs_0 ? 7'h22 : _GEN_2281; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2283 = 10'heb == io_inputs_0 ? 7'h23 : _GEN_2282; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2284 = 10'hec == io_inputs_0 ? 7'h24 : _GEN_2283; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2285 = 10'hed == io_inputs_0 ? 7'h25 : _GEN_2284; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2286 = 10'hee == io_inputs_0 ? 7'h26 : _GEN_2285; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2287 = 10'hef == io_inputs_0 ? 7'h27 : _GEN_2286; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2288 = 10'hf0 == io_inputs_0 ? 7'h28 : _GEN_2287; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2289 = 10'hf1 == io_inputs_0 ? 7'h29 : _GEN_2288; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2290 = 10'hf2 == io_inputs_0 ? 7'h2a : _GEN_2289; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2291 = 10'hf3 == io_inputs_0 ? 7'h2b : _GEN_2290; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2292 = 10'hf4 == io_inputs_0 ? 7'h2c : _GEN_2291; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2293 = 10'hf5 == io_inputs_0 ? 7'h2d : _GEN_2292; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2294 = 10'hf6 == io_inputs_0 ? 7'h2e : _GEN_2293; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2295 = 10'hf7 == io_inputs_0 ? 7'h2f : _GEN_2294; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2296 = 10'hf8 == io_inputs_0 ? 7'h30 : _GEN_2295; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2297 = 10'hf9 == io_inputs_0 ? 7'h31 : _GEN_2296; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2298 = 10'hfa == io_inputs_0 ? 7'h32 : _GEN_2297; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2299 = 10'hfb == io_inputs_0 ? 7'h33 : _GEN_2298; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2300 = 10'hfc == io_inputs_0 ? 7'h34 : _GEN_2299; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2301 = 10'hfd == io_inputs_0 ? 7'h35 : _GEN_2300; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2302 = 10'hfe == io_inputs_0 ? 7'h36 : _GEN_2301; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2303 = 10'hff == io_inputs_0 ? 7'h37 : _GEN_2302; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2304 = 10'h100 == io_inputs_0 ? 7'h38 : _GEN_2303; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2305 = 10'h101 == io_inputs_0 ? 7'h39 : _GEN_2304; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2306 = 10'h102 == io_inputs_0 ? 7'h3a : _GEN_2305; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2307 = 10'h103 == io_inputs_0 ? 7'h3b : _GEN_2306; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2308 = 10'h104 == io_inputs_0 ? 7'h3c : _GEN_2307; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2309 = 10'h105 == io_inputs_0 ? 7'h3d : _GEN_2308; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2310 = 10'h106 == io_inputs_0 ? 7'h3e : _GEN_2309; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2311 = 10'h107 == io_inputs_0 ? 7'h3f : _GEN_2310; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2312 = 10'h108 == io_inputs_0 ? 7'h40 : _GEN_2311; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2313 = 10'h109 == io_inputs_0 ? 7'h41 : _GEN_2312; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2314 = 10'h10a == io_inputs_0 ? 7'h42 : _GEN_2313; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2315 = 10'h10b == io_inputs_0 ? 7'h43 : _GEN_2314; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2316 = 10'h10c == io_inputs_0 ? 7'h44 : _GEN_2315; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2317 = 10'h10d == io_inputs_0 ? 7'h45 : _GEN_2316; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2318 = 10'h10e == io_inputs_0 ? 7'h46 : _GEN_2317; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2319 = 10'h10f == io_inputs_0 ? 7'h47 : _GEN_2318; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2320 = 10'h110 == io_inputs_0 ? 7'h48 : _GEN_2319; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2321 = 10'h111 == io_inputs_0 ? 7'h49 : _GEN_2320; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2322 = 10'h112 == io_inputs_0 ? 7'h4a : _GEN_2321; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2323 = 10'h113 == io_inputs_0 ? 7'h4b : _GEN_2322; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2324 = 10'h114 == io_inputs_0 ? 7'h4c : _GEN_2323; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2325 = 10'h115 == io_inputs_0 ? 7'h4d : _GEN_2324; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2326 = 10'h116 == io_inputs_0 ? 7'h4e : _GEN_2325; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2327 = 10'h117 == io_inputs_0 ? 7'h4f : _GEN_2326; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2328 = 10'h118 == io_inputs_0 ? 7'h50 : _GEN_2327; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2329 = 10'h119 == io_inputs_0 ? 7'h51 : _GEN_2328; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2330 = 10'h11a == io_inputs_0 ? 7'h52 : _GEN_2329; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2331 = 10'h11b == io_inputs_0 ? 7'h53 : _GEN_2330; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2332 = 10'h11c == io_inputs_0 ? 7'h54 : _GEN_2331; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2333 = 10'h11d == io_inputs_0 ? 7'h55 : _GEN_2332; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2334 = 10'h11e == io_inputs_0 ? 7'h56 : _GEN_2333; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2335 = 10'h11f == io_inputs_0 ? 7'h57 : _GEN_2334; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2336 = 10'h120 == io_inputs_0 ? 7'h58 : _GEN_2335; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2337 = 10'h121 == io_inputs_0 ? 7'h59 : _GEN_2336; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2338 = 10'h122 == io_inputs_0 ? 7'h5a : _GEN_2337; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2339 = 10'h123 == io_inputs_0 ? 7'h5b : _GEN_2338; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2340 = 10'h124 == io_inputs_0 ? 7'h5c : _GEN_2339; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2341 = 10'h125 == io_inputs_0 ? 7'h5d : _GEN_2340; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2342 = 10'h126 == io_inputs_0 ? 7'h5e : _GEN_2341; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2343 = 10'h127 == io_inputs_0 ? 7'h5f : _GEN_2342; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2344 = 10'h128 == io_inputs_0 ? 7'h60 : _GEN_2343; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2345 = 10'h129 == io_inputs_0 ? 7'h61 : _GEN_2344; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2346 = 10'h12a == io_inputs_0 ? 7'h62 : _GEN_2345; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2347 = 10'h12b == io_inputs_0 ? 7'h63 : _GEN_2346; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2348 = 10'h12c == io_inputs_0 ? 7'h64 : _GEN_2347; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2349 = 10'h12d == io_inputs_0 ? 7'h0 : _GEN_2348; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2350 = 10'h12e == io_inputs_0 ? 7'h0 : _GEN_2349; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2351 = 10'h12f == io_inputs_0 ? 7'h0 : _GEN_2350; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2352 = 10'h130 == io_inputs_0 ? 7'h0 : _GEN_2351; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2353 = 10'h131 == io_inputs_0 ? 7'h0 : _GEN_2352; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2354 = 10'h132 == io_inputs_0 ? 7'h0 : _GEN_2353; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2355 = 10'h133 == io_inputs_0 ? 7'h0 : _GEN_2354; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2356 = 10'h134 == io_inputs_0 ? 7'h0 : _GEN_2355; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2357 = 10'h135 == io_inputs_0 ? 7'h0 : _GEN_2356; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2358 = 10'h136 == io_inputs_0 ? 7'h0 : _GEN_2357; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2359 = 10'h137 == io_inputs_0 ? 7'h0 : _GEN_2358; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2360 = 10'h138 == io_inputs_0 ? 7'h0 : _GEN_2359; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2361 = 10'h139 == io_inputs_0 ? 7'h0 : _GEN_2360; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2362 = 10'h13a == io_inputs_0 ? 7'h0 : _GEN_2361; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2363 = 10'h13b == io_inputs_0 ? 7'h0 : _GEN_2362; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2364 = 10'h13c == io_inputs_0 ? 7'h0 : _GEN_2363; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2365 = 10'h13d == io_inputs_0 ? 7'h0 : _GEN_2364; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2366 = 10'h13e == io_inputs_0 ? 7'h0 : _GEN_2365; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2367 = 10'h13f == io_inputs_0 ? 7'h0 : _GEN_2366; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2368 = 10'h140 == io_inputs_0 ? 7'h0 : _GEN_2367; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2369 = 10'h141 == io_inputs_0 ? 7'h0 : _GEN_2368; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2370 = 10'h142 == io_inputs_0 ? 7'h0 : _GEN_2369; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2371 = 10'h143 == io_inputs_0 ? 7'h0 : _GEN_2370; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2372 = 10'h144 == io_inputs_0 ? 7'h0 : _GEN_2371; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2373 = 10'h145 == io_inputs_0 ? 7'h0 : _GEN_2372; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2374 = 10'h146 == io_inputs_0 ? 7'h0 : _GEN_2373; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2375 = 10'h147 == io_inputs_0 ? 7'h0 : _GEN_2374; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2376 = 10'h148 == io_inputs_0 ? 7'h0 : _GEN_2375; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2377 = 10'h149 == io_inputs_0 ? 7'h0 : _GEN_2376; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2378 = 10'h14a == io_inputs_0 ? 7'h0 : _GEN_2377; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2379 = 10'h14b == io_inputs_0 ? 7'h0 : _GEN_2378; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2380 = 10'h14c == io_inputs_0 ? 7'h0 : _GEN_2379; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2381 = 10'h14d == io_inputs_0 ? 7'h0 : _GEN_2380; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2382 = 10'h14e == io_inputs_0 ? 7'h0 : _GEN_2381; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2383 = 10'h14f == io_inputs_0 ? 7'h0 : _GEN_2382; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2384 = 10'h150 == io_inputs_0 ? 7'h0 : _GEN_2383; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2385 = 10'h151 == io_inputs_0 ? 7'h0 : _GEN_2384; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2386 = 10'h152 == io_inputs_0 ? 7'h0 : _GEN_2385; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2387 = 10'h153 == io_inputs_0 ? 7'h0 : _GEN_2386; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2388 = 10'h154 == io_inputs_0 ? 7'h0 : _GEN_2387; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2389 = 10'h155 == io_inputs_0 ? 7'h0 : _GEN_2388; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2390 = 10'h156 == io_inputs_0 ? 7'h0 : _GEN_2389; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2391 = 10'h157 == io_inputs_0 ? 7'h0 : _GEN_2390; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2392 = 10'h158 == io_inputs_0 ? 7'h0 : _GEN_2391; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2393 = 10'h159 == io_inputs_0 ? 7'h0 : _GEN_2392; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2394 = 10'h15a == io_inputs_0 ? 7'h0 : _GEN_2393; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2395 = 10'h15b == io_inputs_0 ? 7'h0 : _GEN_2394; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2396 = 10'h15c == io_inputs_0 ? 7'h0 : _GEN_2395; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2397 = 10'h15d == io_inputs_0 ? 7'h0 : _GEN_2396; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2398 = 10'h15e == io_inputs_0 ? 7'h0 : _GEN_2397; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2399 = 10'h15f == io_inputs_0 ? 7'h0 : _GEN_2398; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2400 = 10'h160 == io_inputs_0 ? 7'h0 : _GEN_2399; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2401 = 10'h161 == io_inputs_0 ? 7'h0 : _GEN_2400; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2402 = 10'h162 == io_inputs_0 ? 7'h0 : _GEN_2401; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2403 = 10'h163 == io_inputs_0 ? 7'h0 : _GEN_2402; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2404 = 10'h164 == io_inputs_0 ? 7'h0 : _GEN_2403; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2405 = 10'h165 == io_inputs_0 ? 7'h0 : _GEN_2404; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2406 = 10'h166 == io_inputs_0 ? 7'h0 : _GEN_2405; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2407 = 10'h167 == io_inputs_0 ? 7'h0 : _GEN_2406; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2408 = 10'h168 == io_inputs_0 ? 7'h0 : _GEN_2407; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2409 = 10'h169 == io_inputs_0 ? 7'h0 : _GEN_2408; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2410 = 10'h16a == io_inputs_0 ? 7'h0 : _GEN_2409; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2411 = 10'h16b == io_inputs_0 ? 7'h0 : _GEN_2410; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2412 = 10'h16c == io_inputs_0 ? 7'h0 : _GEN_2411; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2413 = 10'h16d == io_inputs_0 ? 7'h0 : _GEN_2412; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2414 = 10'h16e == io_inputs_0 ? 7'h0 : _GEN_2413; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2415 = 10'h16f == io_inputs_0 ? 7'h0 : _GEN_2414; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2416 = 10'h170 == io_inputs_0 ? 7'h0 : _GEN_2415; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2417 = 10'h171 == io_inputs_0 ? 7'h0 : _GEN_2416; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2418 = 10'h172 == io_inputs_0 ? 7'h0 : _GEN_2417; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2419 = 10'h173 == io_inputs_0 ? 7'h0 : _GEN_2418; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2420 = 10'h174 == io_inputs_0 ? 7'h0 : _GEN_2419; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2421 = 10'h175 == io_inputs_0 ? 7'h0 : _GEN_2420; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2422 = 10'h176 == io_inputs_0 ? 7'h0 : _GEN_2421; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2423 = 10'h177 == io_inputs_0 ? 7'h0 : _GEN_2422; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2424 = 10'h178 == io_inputs_0 ? 7'h0 : _GEN_2423; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2425 = 10'h179 == io_inputs_0 ? 7'h0 : _GEN_2424; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2426 = 10'h17a == io_inputs_0 ? 7'h0 : _GEN_2425; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2427 = 10'h17b == io_inputs_0 ? 7'h0 : _GEN_2426; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2428 = 10'h17c == io_inputs_0 ? 7'h0 : _GEN_2427; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2429 = 10'h17d == io_inputs_0 ? 7'h0 : _GEN_2428; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2430 = 10'h17e == io_inputs_0 ? 7'h0 : _GEN_2429; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2431 = 10'h17f == io_inputs_0 ? 7'h0 : _GEN_2430; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2432 = 10'h180 == io_inputs_0 ? 7'h0 : _GEN_2431; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2433 = 10'h181 == io_inputs_0 ? 7'h0 : _GEN_2432; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2434 = 10'h182 == io_inputs_0 ? 7'h0 : _GEN_2433; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2435 = 10'h183 == io_inputs_0 ? 7'h0 : _GEN_2434; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2436 = 10'h184 == io_inputs_0 ? 7'h0 : _GEN_2435; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2437 = 10'h185 == io_inputs_0 ? 7'h0 : _GEN_2436; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2438 = 10'h186 == io_inputs_0 ? 7'h0 : _GEN_2437; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2439 = 10'h187 == io_inputs_0 ? 7'h0 : _GEN_2438; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2440 = 10'h188 == io_inputs_0 ? 7'h0 : _GEN_2439; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2441 = 10'h189 == io_inputs_0 ? 7'h0 : _GEN_2440; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2442 = 10'h18a == io_inputs_0 ? 7'h0 : _GEN_2441; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2443 = 10'h18b == io_inputs_0 ? 7'h0 : _GEN_2442; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2444 = 10'h18c == io_inputs_0 ? 7'h0 : _GEN_2443; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2445 = 10'h18d == io_inputs_0 ? 7'h0 : _GEN_2444; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2446 = 10'h18e == io_inputs_0 ? 7'h0 : _GEN_2445; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2447 = 10'h18f == io_inputs_0 ? 7'h0 : _GEN_2446; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2448 = 10'h190 == io_inputs_0 ? 7'h0 : _GEN_2447; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2449 = 10'h191 == io_inputs_0 ? 7'h0 : _GEN_2448; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2450 = 10'h192 == io_inputs_0 ? 7'h0 : _GEN_2449; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2451 = 10'h193 == io_inputs_0 ? 7'h0 : _GEN_2450; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2452 = 10'h194 == io_inputs_0 ? 7'h0 : _GEN_2451; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2453 = 10'h195 == io_inputs_0 ? 7'h0 : _GEN_2452; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2454 = 10'h196 == io_inputs_0 ? 7'h0 : _GEN_2453; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2455 = 10'h197 == io_inputs_0 ? 7'h0 : _GEN_2454; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2456 = 10'h198 == io_inputs_0 ? 7'h0 : _GEN_2455; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2457 = 10'h199 == io_inputs_0 ? 7'h0 : _GEN_2456; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2458 = 10'h19a == io_inputs_0 ? 7'h0 : _GEN_2457; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2459 = 10'h19b == io_inputs_0 ? 7'h0 : _GEN_2458; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2460 = 10'h19c == io_inputs_0 ? 7'h0 : _GEN_2459; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2461 = 10'h19d == io_inputs_0 ? 7'h0 : _GEN_2460; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2462 = 10'h19e == io_inputs_0 ? 7'h0 : _GEN_2461; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2463 = 10'h19f == io_inputs_0 ? 7'h0 : _GEN_2462; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2464 = 10'h1a0 == io_inputs_0 ? 7'h0 : _GEN_2463; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2465 = 10'h1a1 == io_inputs_0 ? 7'h0 : _GEN_2464; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2466 = 10'h1a2 == io_inputs_0 ? 7'h0 : _GEN_2465; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2467 = 10'h1a3 == io_inputs_0 ? 7'h0 : _GEN_2466; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2468 = 10'h1a4 == io_inputs_0 ? 7'h0 : _GEN_2467; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2469 = 10'h1a5 == io_inputs_0 ? 7'h0 : _GEN_2468; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2470 = 10'h1a6 == io_inputs_0 ? 7'h0 : _GEN_2469; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2471 = 10'h1a7 == io_inputs_0 ? 7'h0 : _GEN_2470; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2472 = 10'h1a8 == io_inputs_0 ? 7'h0 : _GEN_2471; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2473 = 10'h1a9 == io_inputs_0 ? 7'h0 : _GEN_2472; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2474 = 10'h1aa == io_inputs_0 ? 7'h0 : _GEN_2473; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2475 = 10'h1ab == io_inputs_0 ? 7'h0 : _GEN_2474; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2476 = 10'h1ac == io_inputs_0 ? 7'h0 : _GEN_2475; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2477 = 10'h1ad == io_inputs_0 ? 7'h0 : _GEN_2476; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2478 = 10'h1ae == io_inputs_0 ? 7'h0 : _GEN_2477; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2479 = 10'h1af == io_inputs_0 ? 7'h0 : _GEN_2478; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2480 = 10'h1b0 == io_inputs_0 ? 7'h0 : _GEN_2479; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2481 = 10'h1b1 == io_inputs_0 ? 7'h0 : _GEN_2480; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2482 = 10'h1b2 == io_inputs_0 ? 7'h0 : _GEN_2481; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2483 = 10'h1b3 == io_inputs_0 ? 7'h0 : _GEN_2482; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2484 = 10'h1b4 == io_inputs_0 ? 7'h0 : _GEN_2483; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2485 = 10'h1b5 == io_inputs_0 ? 7'h0 : _GEN_2484; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2486 = 10'h1b6 == io_inputs_0 ? 7'h0 : _GEN_2485; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2487 = 10'h1b7 == io_inputs_0 ? 7'h0 : _GEN_2486; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2488 = 10'h1b8 == io_inputs_0 ? 7'h0 : _GEN_2487; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2489 = 10'h1b9 == io_inputs_0 ? 7'h0 : _GEN_2488; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2490 = 10'h1ba == io_inputs_0 ? 7'h0 : _GEN_2489; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2491 = 10'h1bb == io_inputs_0 ? 7'h0 : _GEN_2490; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2492 = 10'h1bc == io_inputs_0 ? 7'h0 : _GEN_2491; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2493 = 10'h1bd == io_inputs_0 ? 7'h0 : _GEN_2492; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2494 = 10'h1be == io_inputs_0 ? 7'h0 : _GEN_2493; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2495 = 10'h1bf == io_inputs_0 ? 7'h0 : _GEN_2494; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2496 = 10'h1c0 == io_inputs_0 ? 7'h0 : _GEN_2495; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2497 = 10'h1c1 == io_inputs_0 ? 7'h0 : _GEN_2496; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2498 = 10'h1c2 == io_inputs_0 ? 7'h0 : _GEN_2497; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2499 = 10'h1c3 == io_inputs_0 ? 7'h0 : _GEN_2498; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2500 = 10'h1c4 == io_inputs_0 ? 7'h0 : _GEN_2499; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2501 = 10'h1c5 == io_inputs_0 ? 7'h0 : _GEN_2500; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2502 = 10'h1c6 == io_inputs_0 ? 7'h0 : _GEN_2501; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2503 = 10'h1c7 == io_inputs_0 ? 7'h0 : _GEN_2502; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2504 = 10'h1c8 == io_inputs_0 ? 7'h0 : _GEN_2503; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2505 = 10'h1c9 == io_inputs_0 ? 7'h0 : _GEN_2504; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2506 = 10'h1ca == io_inputs_0 ? 7'h0 : _GEN_2505; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2507 = 10'h1cb == io_inputs_0 ? 7'h0 : _GEN_2506; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2508 = 10'h1cc == io_inputs_0 ? 7'h0 : _GEN_2507; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2509 = 10'h1cd == io_inputs_0 ? 7'h0 : _GEN_2508; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2510 = 10'h1ce == io_inputs_0 ? 7'h0 : _GEN_2509; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2511 = 10'h1cf == io_inputs_0 ? 7'h0 : _GEN_2510; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2512 = 10'h1d0 == io_inputs_0 ? 7'h0 : _GEN_2511; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2513 = 10'h1d1 == io_inputs_0 ? 7'h0 : _GEN_2512; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2514 = 10'h1d2 == io_inputs_0 ? 7'h0 : _GEN_2513; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2515 = 10'h1d3 == io_inputs_0 ? 7'h0 : _GEN_2514; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2516 = 10'h1d4 == io_inputs_0 ? 7'h0 : _GEN_2515; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2517 = 10'h1d5 == io_inputs_0 ? 7'h0 : _GEN_2516; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2518 = 10'h1d6 == io_inputs_0 ? 7'h0 : _GEN_2517; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2519 = 10'h1d7 == io_inputs_0 ? 7'h0 : _GEN_2518; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2520 = 10'h1d8 == io_inputs_0 ? 7'h0 : _GEN_2519; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2521 = 10'h1d9 == io_inputs_0 ? 7'h0 : _GEN_2520; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2522 = 10'h1da == io_inputs_0 ? 7'h0 : _GEN_2521; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2523 = 10'h1db == io_inputs_0 ? 7'h0 : _GEN_2522; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2524 = 10'h1dc == io_inputs_0 ? 7'h0 : _GEN_2523; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2525 = 10'h1dd == io_inputs_0 ? 7'h0 : _GEN_2524; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2526 = 10'h1de == io_inputs_0 ? 7'h0 : _GEN_2525; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2527 = 10'h1df == io_inputs_0 ? 7'h0 : _GEN_2526; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2528 = 10'h1e0 == io_inputs_0 ? 7'h0 : _GEN_2527; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2529 = 10'h1e1 == io_inputs_0 ? 7'h0 : _GEN_2528; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2530 = 10'h1e2 == io_inputs_0 ? 7'h0 : _GEN_2529; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2531 = 10'h1e3 == io_inputs_0 ? 7'h0 : _GEN_2530; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2532 = 10'h1e4 == io_inputs_0 ? 7'h0 : _GEN_2531; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2533 = 10'h1e5 == io_inputs_0 ? 7'h0 : _GEN_2532; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2534 = 10'h1e6 == io_inputs_0 ? 7'h0 : _GEN_2533; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2535 = 10'h1e7 == io_inputs_0 ? 7'h0 : _GEN_2534; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2536 = 10'h1e8 == io_inputs_0 ? 7'h0 : _GEN_2535; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2537 = 10'h1e9 == io_inputs_0 ? 7'h0 : _GEN_2536; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2538 = 10'h1ea == io_inputs_0 ? 7'h0 : _GEN_2537; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2539 = 10'h1eb == io_inputs_0 ? 7'h0 : _GEN_2538; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2540 = 10'h1ec == io_inputs_0 ? 7'h0 : _GEN_2539; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2541 = 10'h1ed == io_inputs_0 ? 7'h0 : _GEN_2540; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2542 = 10'h1ee == io_inputs_0 ? 7'h0 : _GEN_2541; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2543 = 10'h1ef == io_inputs_0 ? 7'h0 : _GEN_2542; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2544 = 10'h1f0 == io_inputs_0 ? 7'h0 : _GEN_2543; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2545 = 10'h1f1 == io_inputs_0 ? 7'h0 : _GEN_2544; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2546 = 10'h1f2 == io_inputs_0 ? 7'h0 : _GEN_2545; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2547 = 10'h1f3 == io_inputs_0 ? 7'h0 : _GEN_2546; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2548 = 10'h1f4 == io_inputs_0 ? 7'h0 : _GEN_2547; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2549 = 10'h1f5 == io_inputs_0 ? 7'h0 : _GEN_2548; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2550 = 10'h1f6 == io_inputs_0 ? 7'h0 : _GEN_2549; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2551 = 10'h1f7 == io_inputs_0 ? 7'h0 : _GEN_2550; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2552 = 10'h1f8 == io_inputs_0 ? 7'h0 : _GEN_2551; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2553 = 10'h1f9 == io_inputs_0 ? 7'h0 : _GEN_2552; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2554 = 10'h1fa == io_inputs_0 ? 7'h0 : _GEN_2553; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2555 = 10'h1fb == io_inputs_0 ? 7'h0 : _GEN_2554; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2556 = 10'h1fc == io_inputs_0 ? 7'h0 : _GEN_2555; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2557 = 10'h1fd == io_inputs_0 ? 7'h0 : _GEN_2556; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2558 = 10'h1fe == io_inputs_0 ? 7'h0 : _GEN_2557; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2559 = 10'h1ff == io_inputs_0 ? 7'h0 : _GEN_2558; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2560 = 10'h200 == io_inputs_0 ? 7'h0 : _GEN_2559; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2561 = 10'h201 == io_inputs_0 ? 7'h0 : _GEN_2560; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2562 = 10'h202 == io_inputs_0 ? 7'h0 : _GEN_2561; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2563 = 10'h203 == io_inputs_0 ? 7'h0 : _GEN_2562; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2564 = 10'h204 == io_inputs_0 ? 7'h0 : _GEN_2563; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2565 = 10'h205 == io_inputs_0 ? 7'h0 : _GEN_2564; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2566 = 10'h206 == io_inputs_0 ? 7'h0 : _GEN_2565; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2567 = 10'h207 == io_inputs_0 ? 7'h0 : _GEN_2566; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2568 = 10'h208 == io_inputs_0 ? 7'h0 : _GEN_2567; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2569 = 10'h209 == io_inputs_0 ? 7'h0 : _GEN_2568; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2570 = 10'h20a == io_inputs_0 ? 7'h0 : _GEN_2569; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2571 = 10'h20b == io_inputs_0 ? 7'h0 : _GEN_2570; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2572 = 10'h20c == io_inputs_0 ? 7'h0 : _GEN_2571; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2573 = 10'h20d == io_inputs_0 ? 7'h0 : _GEN_2572; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2574 = 10'h20e == io_inputs_0 ? 7'h0 : _GEN_2573; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2575 = 10'h20f == io_inputs_0 ? 7'h0 : _GEN_2574; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2576 = 10'h210 == io_inputs_0 ? 7'h0 : _GEN_2575; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2577 = 10'h211 == io_inputs_0 ? 7'h0 : _GEN_2576; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2578 = 10'h212 == io_inputs_0 ? 7'h0 : _GEN_2577; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2579 = 10'h213 == io_inputs_0 ? 7'h0 : _GEN_2578; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2580 = 10'h214 == io_inputs_0 ? 7'h0 : _GEN_2579; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2581 = 10'h215 == io_inputs_0 ? 7'h0 : _GEN_2580; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2582 = 10'h216 == io_inputs_0 ? 7'h0 : _GEN_2581; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2583 = 10'h217 == io_inputs_0 ? 7'h0 : _GEN_2582; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2584 = 10'h218 == io_inputs_0 ? 7'h0 : _GEN_2583; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2585 = 10'h219 == io_inputs_0 ? 7'h0 : _GEN_2584; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2586 = 10'h21a == io_inputs_0 ? 7'h0 : _GEN_2585; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2587 = 10'h21b == io_inputs_0 ? 7'h0 : _GEN_2586; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2588 = 10'h21c == io_inputs_0 ? 7'h0 : _GEN_2587; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2589 = 10'h21d == io_inputs_0 ? 7'h0 : _GEN_2588; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2590 = 10'h21e == io_inputs_0 ? 7'h0 : _GEN_2589; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2591 = 10'h21f == io_inputs_0 ? 7'h0 : _GEN_2590; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2592 = 10'h220 == io_inputs_0 ? 7'h0 : _GEN_2591; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2593 = 10'h221 == io_inputs_0 ? 7'h0 : _GEN_2592; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2594 = 10'h222 == io_inputs_0 ? 7'h0 : _GEN_2593; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2595 = 10'h223 == io_inputs_0 ? 7'h0 : _GEN_2594; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2596 = 10'h224 == io_inputs_0 ? 7'h0 : _GEN_2595; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2597 = 10'h225 == io_inputs_0 ? 7'h0 : _GEN_2596; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2598 = 10'h226 == io_inputs_0 ? 7'h0 : _GEN_2597; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2599 = 10'h227 == io_inputs_0 ? 7'h0 : _GEN_2598; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2600 = 10'h228 == io_inputs_0 ? 7'h0 : _GEN_2599; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2601 = 10'h229 == io_inputs_0 ? 7'h0 : _GEN_2600; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2602 = 10'h22a == io_inputs_0 ? 7'h0 : _GEN_2601; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2603 = 10'h22b == io_inputs_0 ? 7'h0 : _GEN_2602; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2604 = 10'h22c == io_inputs_0 ? 7'h0 : _GEN_2603; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2605 = 10'h22d == io_inputs_0 ? 7'h0 : _GEN_2604; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2606 = 10'h22e == io_inputs_0 ? 7'h0 : _GEN_2605; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2607 = 10'h22f == io_inputs_0 ? 7'h0 : _GEN_2606; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2608 = 10'h230 == io_inputs_0 ? 7'h0 : _GEN_2607; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2609 = 10'h231 == io_inputs_0 ? 7'h0 : _GEN_2608; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2610 = 10'h232 == io_inputs_0 ? 7'h0 : _GEN_2609; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2611 = 10'h233 == io_inputs_0 ? 7'h0 : _GEN_2610; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2612 = 10'h234 == io_inputs_0 ? 7'h0 : _GEN_2611; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2613 = 10'h235 == io_inputs_0 ? 7'h0 : _GEN_2612; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2614 = 10'h236 == io_inputs_0 ? 7'h0 : _GEN_2613; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2615 = 10'h237 == io_inputs_0 ? 7'h0 : _GEN_2614; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2616 = 10'h238 == io_inputs_0 ? 7'h0 : _GEN_2615; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2617 = 10'h239 == io_inputs_0 ? 7'h0 : _GEN_2616; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2618 = 10'h23a == io_inputs_0 ? 7'h0 : _GEN_2617; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2619 = 10'h23b == io_inputs_0 ? 7'h0 : _GEN_2618; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2620 = 10'h23c == io_inputs_0 ? 7'h0 : _GEN_2619; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2621 = 10'h23d == io_inputs_0 ? 7'h0 : _GEN_2620; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2622 = 10'h23e == io_inputs_0 ? 7'h0 : _GEN_2621; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2623 = 10'h23f == io_inputs_0 ? 7'h0 : _GEN_2622; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2624 = 10'h240 == io_inputs_0 ? 7'h0 : _GEN_2623; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2625 = 10'h241 == io_inputs_0 ? 7'h0 : _GEN_2624; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2626 = 10'h242 == io_inputs_0 ? 7'h0 : _GEN_2625; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2627 = 10'h243 == io_inputs_0 ? 7'h0 : _GEN_2626; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2628 = 10'h244 == io_inputs_0 ? 7'h0 : _GEN_2627; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2629 = 10'h245 == io_inputs_0 ? 7'h0 : _GEN_2628; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2630 = 10'h246 == io_inputs_0 ? 7'h0 : _GEN_2629; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2631 = 10'h247 == io_inputs_0 ? 7'h0 : _GEN_2630; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2632 = 10'h248 == io_inputs_0 ? 7'h0 : _GEN_2631; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2633 = 10'h249 == io_inputs_0 ? 7'h0 : _GEN_2632; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2634 = 10'h24a == io_inputs_0 ? 7'h0 : _GEN_2633; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2635 = 10'h24b == io_inputs_0 ? 7'h0 : _GEN_2634; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2636 = 10'h24c == io_inputs_0 ? 7'h0 : _GEN_2635; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2637 = 10'h24d == io_inputs_0 ? 7'h0 : _GEN_2636; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2638 = 10'h24e == io_inputs_0 ? 7'h0 : _GEN_2637; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2639 = 10'h24f == io_inputs_0 ? 7'h0 : _GEN_2638; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2640 = 10'h250 == io_inputs_0 ? 7'h0 : _GEN_2639; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2641 = 10'h251 == io_inputs_0 ? 7'h0 : _GEN_2640; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2642 = 10'h252 == io_inputs_0 ? 7'h0 : _GEN_2641; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2643 = 10'h253 == io_inputs_0 ? 7'h0 : _GEN_2642; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2644 = 10'h254 == io_inputs_0 ? 7'h0 : _GEN_2643; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2645 = 10'h255 == io_inputs_0 ? 7'h0 : _GEN_2644; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2646 = 10'h256 == io_inputs_0 ? 7'h0 : _GEN_2645; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2647 = 10'h257 == io_inputs_0 ? 7'h0 : _GEN_2646; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2648 = 10'h258 == io_inputs_0 ? 7'h0 : _GEN_2647; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2649 = 10'h259 == io_inputs_0 ? 7'h0 : _GEN_2648; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2650 = 10'h25a == io_inputs_0 ? 7'h0 : _GEN_2649; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2651 = 10'h25b == io_inputs_0 ? 7'h0 : _GEN_2650; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2652 = 10'h25c == io_inputs_0 ? 7'h0 : _GEN_2651; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2653 = 10'h25d == io_inputs_0 ? 7'h0 : _GEN_2652; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2654 = 10'h25e == io_inputs_0 ? 7'h0 : _GEN_2653; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2655 = 10'h25f == io_inputs_0 ? 7'h0 : _GEN_2654; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2656 = 10'h260 == io_inputs_0 ? 7'h0 : _GEN_2655; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2657 = 10'h261 == io_inputs_0 ? 7'h0 : _GEN_2656; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2658 = 10'h262 == io_inputs_0 ? 7'h0 : _GEN_2657; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2659 = 10'h263 == io_inputs_0 ? 7'h0 : _GEN_2658; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2660 = 10'h264 == io_inputs_0 ? 7'h0 : _GEN_2659; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2661 = 10'h265 == io_inputs_0 ? 7'h0 : _GEN_2660; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2662 = 10'h266 == io_inputs_0 ? 7'h0 : _GEN_2661; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2663 = 10'h267 == io_inputs_0 ? 7'h0 : _GEN_2662; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2664 = 10'h268 == io_inputs_0 ? 7'h0 : _GEN_2663; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2665 = 10'h269 == io_inputs_0 ? 7'h0 : _GEN_2664; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2666 = 10'h26a == io_inputs_0 ? 7'h0 : _GEN_2665; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2667 = 10'h26b == io_inputs_0 ? 7'h0 : _GEN_2666; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2668 = 10'h26c == io_inputs_0 ? 7'h0 : _GEN_2667; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2669 = 10'h26d == io_inputs_0 ? 7'h0 : _GEN_2668; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2670 = 10'h26e == io_inputs_0 ? 7'h0 : _GEN_2669; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2671 = 10'h26f == io_inputs_0 ? 7'h0 : _GEN_2670; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2672 = 10'h270 == io_inputs_0 ? 7'h0 : _GEN_2671; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2673 = 10'h271 == io_inputs_0 ? 7'h0 : _GEN_2672; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2674 = 10'h272 == io_inputs_0 ? 7'h0 : _GEN_2673; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2675 = 10'h273 == io_inputs_0 ? 7'h0 : _GEN_2674; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2676 = 10'h274 == io_inputs_0 ? 7'h0 : _GEN_2675; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2677 = 10'h275 == io_inputs_0 ? 7'h0 : _GEN_2676; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2678 = 10'h276 == io_inputs_0 ? 7'h0 : _GEN_2677; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2679 = 10'h277 == io_inputs_0 ? 7'h0 : _GEN_2678; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2680 = 10'h278 == io_inputs_0 ? 7'h0 : _GEN_2679; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2681 = 10'h279 == io_inputs_0 ? 7'h0 : _GEN_2680; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2682 = 10'h27a == io_inputs_0 ? 7'h0 : _GEN_2681; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2683 = 10'h27b == io_inputs_0 ? 7'h0 : _GEN_2682; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2684 = 10'h27c == io_inputs_0 ? 7'h0 : _GEN_2683; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2685 = 10'h27d == io_inputs_0 ? 7'h0 : _GEN_2684; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2686 = 10'h27e == io_inputs_0 ? 7'h0 : _GEN_2685; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2687 = 10'h27f == io_inputs_0 ? 7'h0 : _GEN_2686; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2688 = 10'h280 == io_inputs_0 ? 7'h0 : _GEN_2687; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2689 = 10'h281 == io_inputs_0 ? 7'h0 : _GEN_2688; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2690 = 10'h282 == io_inputs_0 ? 7'h0 : _GEN_2689; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2691 = 10'h283 == io_inputs_0 ? 7'h0 : _GEN_2690; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2692 = 10'h284 == io_inputs_0 ? 7'h0 : _GEN_2691; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2693 = 10'h285 == io_inputs_0 ? 7'h0 : _GEN_2692; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2694 = 10'h286 == io_inputs_0 ? 7'h0 : _GEN_2693; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2695 = 10'h287 == io_inputs_0 ? 7'h0 : _GEN_2694; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2696 = 10'h288 == io_inputs_0 ? 7'h0 : _GEN_2695; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2697 = 10'h289 == io_inputs_0 ? 7'h0 : _GEN_2696; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2698 = 10'h28a == io_inputs_0 ? 7'h0 : _GEN_2697; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2699 = 10'h28b == io_inputs_0 ? 7'h0 : _GEN_2698; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2700 = 10'h28c == io_inputs_0 ? 7'h0 : _GEN_2699; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2701 = 10'h28d == io_inputs_0 ? 7'h0 : _GEN_2700; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2702 = 10'h28e == io_inputs_0 ? 7'h0 : _GEN_2701; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2703 = 10'h28f == io_inputs_0 ? 7'h0 : _GEN_2702; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2704 = 10'h290 == io_inputs_0 ? 7'h0 : _GEN_2703; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2705 = 10'h291 == io_inputs_0 ? 7'h0 : _GEN_2704; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2706 = 10'h292 == io_inputs_0 ? 7'h0 : _GEN_2705; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2707 = 10'h293 == io_inputs_0 ? 7'h0 : _GEN_2706; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2708 = 10'h294 == io_inputs_0 ? 7'h0 : _GEN_2707; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2709 = 10'h295 == io_inputs_0 ? 7'h0 : _GEN_2708; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2710 = 10'h296 == io_inputs_0 ? 7'h0 : _GEN_2709; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2711 = 10'h297 == io_inputs_0 ? 7'h0 : _GEN_2710; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2712 = 10'h298 == io_inputs_0 ? 7'h0 : _GEN_2711; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2713 = 10'h299 == io_inputs_0 ? 7'h0 : _GEN_2712; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2714 = 10'h29a == io_inputs_0 ? 7'h0 : _GEN_2713; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2715 = 10'h29b == io_inputs_0 ? 7'h0 : _GEN_2714; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2716 = 10'h29c == io_inputs_0 ? 7'h0 : _GEN_2715; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2717 = 10'h29d == io_inputs_0 ? 7'h0 : _GEN_2716; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2718 = 10'h29e == io_inputs_0 ? 7'h0 : _GEN_2717; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2719 = 10'h29f == io_inputs_0 ? 7'h0 : _GEN_2718; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2720 = 10'h2a0 == io_inputs_0 ? 7'h0 : _GEN_2719; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2721 = 10'h2a1 == io_inputs_0 ? 7'h0 : _GEN_2720; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2722 = 10'h2a2 == io_inputs_0 ? 7'h0 : _GEN_2721; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2723 = 10'h2a3 == io_inputs_0 ? 7'h0 : _GEN_2722; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2724 = 10'h2a4 == io_inputs_0 ? 7'h0 : _GEN_2723; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2725 = 10'h2a5 == io_inputs_0 ? 7'h0 : _GEN_2724; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2726 = 10'h2a6 == io_inputs_0 ? 7'h0 : _GEN_2725; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2727 = 10'h2a7 == io_inputs_0 ? 7'h0 : _GEN_2726; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2728 = 10'h2a8 == io_inputs_0 ? 7'h0 : _GEN_2727; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2729 = 10'h2a9 == io_inputs_0 ? 7'h0 : _GEN_2728; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2730 = 10'h2aa == io_inputs_0 ? 7'h0 : _GEN_2729; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2731 = 10'h2ab == io_inputs_0 ? 7'h0 : _GEN_2730; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2732 = 10'h2ac == io_inputs_0 ? 7'h0 : _GEN_2731; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2733 = 10'h2ad == io_inputs_0 ? 7'h0 : _GEN_2732; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2734 = 10'h2ae == io_inputs_0 ? 7'h0 : _GEN_2733; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2735 = 10'h2af == io_inputs_0 ? 7'h0 : _GEN_2734; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2736 = 10'h2b0 == io_inputs_0 ? 7'h0 : _GEN_2735; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2737 = 10'h2b1 == io_inputs_0 ? 7'h0 : _GEN_2736; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2738 = 10'h2b2 == io_inputs_0 ? 7'h0 : _GEN_2737; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2739 = 10'h2b3 == io_inputs_0 ? 7'h0 : _GEN_2738; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2740 = 10'h2b4 == io_inputs_0 ? 7'h0 : _GEN_2739; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2741 = 10'h2b5 == io_inputs_0 ? 7'h0 : _GEN_2740; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2742 = 10'h2b6 == io_inputs_0 ? 7'h0 : _GEN_2741; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2743 = 10'h2b7 == io_inputs_0 ? 7'h0 : _GEN_2742; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2744 = 10'h2b8 == io_inputs_0 ? 7'h0 : _GEN_2743; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2745 = 10'h2b9 == io_inputs_0 ? 7'h0 : _GEN_2744; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2746 = 10'h2ba == io_inputs_0 ? 7'h0 : _GEN_2745; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2747 = 10'h2bb == io_inputs_0 ? 7'h0 : _GEN_2746; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2748 = 10'h2bc == io_inputs_0 ? 7'h0 : _GEN_2747; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2749 = 10'h2bd == io_inputs_0 ? 7'h0 : _GEN_2748; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2750 = 10'h2be == io_inputs_0 ? 7'h0 : _GEN_2749; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2751 = 10'h2bf == io_inputs_0 ? 7'h0 : _GEN_2750; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2752 = 10'h2c0 == io_inputs_0 ? 7'h0 : _GEN_2751; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2753 = 10'h2c1 == io_inputs_0 ? 7'h0 : _GEN_2752; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2754 = 10'h2c2 == io_inputs_0 ? 7'h0 : _GEN_2753; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2755 = 10'h2c3 == io_inputs_0 ? 7'h0 : _GEN_2754; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2756 = 10'h2c4 == io_inputs_0 ? 7'h0 : _GEN_2755; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2757 = 10'h2c5 == io_inputs_0 ? 7'h0 : _GEN_2756; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2758 = 10'h2c6 == io_inputs_0 ? 7'h0 : _GEN_2757; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2759 = 10'h2c7 == io_inputs_0 ? 7'h0 : _GEN_2758; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2760 = 10'h2c8 == io_inputs_0 ? 7'h0 : _GEN_2759; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2761 = 10'h2c9 == io_inputs_0 ? 7'h0 : _GEN_2760; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2762 = 10'h2ca == io_inputs_0 ? 7'h0 : _GEN_2761; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2763 = 10'h2cb == io_inputs_0 ? 7'h0 : _GEN_2762; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2764 = 10'h2cc == io_inputs_0 ? 7'h0 : _GEN_2763; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2765 = 10'h2cd == io_inputs_0 ? 7'h0 : _GEN_2764; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2766 = 10'h2ce == io_inputs_0 ? 7'h0 : _GEN_2765; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2767 = 10'h2cf == io_inputs_0 ? 7'h0 : _GEN_2766; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2768 = 10'h2d0 == io_inputs_0 ? 7'h0 : _GEN_2767; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2769 = 10'h2d1 == io_inputs_0 ? 7'h0 : _GEN_2768; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2770 = 10'h2d2 == io_inputs_0 ? 7'h0 : _GEN_2769; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2771 = 10'h2d3 == io_inputs_0 ? 7'h0 : _GEN_2770; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2772 = 10'h2d4 == io_inputs_0 ? 7'h0 : _GEN_2771; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2773 = 10'h2d5 == io_inputs_0 ? 7'h0 : _GEN_2772; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2774 = 10'h2d6 == io_inputs_0 ? 7'h0 : _GEN_2773; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2775 = 10'h2d7 == io_inputs_0 ? 7'h0 : _GEN_2774; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2776 = 10'h2d8 == io_inputs_0 ? 7'h0 : _GEN_2775; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2777 = 10'h2d9 == io_inputs_0 ? 7'h0 : _GEN_2776; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2778 = 10'h2da == io_inputs_0 ? 7'h0 : _GEN_2777; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2779 = 10'h2db == io_inputs_0 ? 7'h0 : _GEN_2778; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2780 = 10'h2dc == io_inputs_0 ? 7'h0 : _GEN_2779; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2781 = 10'h2dd == io_inputs_0 ? 7'h0 : _GEN_2780; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2782 = 10'h2de == io_inputs_0 ? 7'h0 : _GEN_2781; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2783 = 10'h2df == io_inputs_0 ? 7'h0 : _GEN_2782; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2784 = 10'h2e0 == io_inputs_0 ? 7'h0 : _GEN_2783; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2785 = 10'h2e1 == io_inputs_0 ? 7'h0 : _GEN_2784; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2786 = 10'h2e2 == io_inputs_0 ? 7'h0 : _GEN_2785; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2787 = 10'h2e3 == io_inputs_0 ? 7'h0 : _GEN_2786; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2788 = 10'h2e4 == io_inputs_0 ? 7'h0 : _GEN_2787; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2789 = 10'h2e5 == io_inputs_0 ? 7'h0 : _GEN_2788; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2790 = 10'h2e6 == io_inputs_0 ? 7'h0 : _GEN_2789; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2791 = 10'h2e7 == io_inputs_0 ? 7'h0 : _GEN_2790; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2792 = 10'h2e8 == io_inputs_0 ? 7'h0 : _GEN_2791; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2793 = 10'h2e9 == io_inputs_0 ? 7'h0 : _GEN_2792; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2794 = 10'h2ea == io_inputs_0 ? 7'h0 : _GEN_2793; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2795 = 10'h2eb == io_inputs_0 ? 7'h0 : _GEN_2794; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2796 = 10'h2ec == io_inputs_0 ? 7'h0 : _GEN_2795; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2797 = 10'h2ed == io_inputs_0 ? 7'h0 : _GEN_2796; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2798 = 10'h2ee == io_inputs_0 ? 7'h0 : _GEN_2797; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2799 = 10'h2ef == io_inputs_0 ? 7'h0 : _GEN_2798; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2800 = 10'h2f0 == io_inputs_0 ? 7'h0 : _GEN_2799; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2801 = 10'h2f1 == io_inputs_0 ? 7'h0 : _GEN_2800; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2802 = 10'h2f2 == io_inputs_0 ? 7'h0 : _GEN_2801; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2803 = 10'h2f3 == io_inputs_0 ? 7'h0 : _GEN_2802; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2804 = 10'h2f4 == io_inputs_0 ? 7'h0 : _GEN_2803; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2805 = 10'h2f5 == io_inputs_0 ? 7'h0 : _GEN_2804; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2806 = 10'h2f6 == io_inputs_0 ? 7'h0 : _GEN_2805; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2807 = 10'h2f7 == io_inputs_0 ? 7'h0 : _GEN_2806; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2808 = 10'h2f8 == io_inputs_0 ? 7'h0 : _GEN_2807; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2809 = 10'h2f9 == io_inputs_0 ? 7'h0 : _GEN_2808; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2810 = 10'h2fa == io_inputs_0 ? 7'h0 : _GEN_2809; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2811 = 10'h2fb == io_inputs_0 ? 7'h0 : _GEN_2810; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2812 = 10'h2fc == io_inputs_0 ? 7'h0 : _GEN_2811; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2813 = 10'h2fd == io_inputs_0 ? 7'h0 : _GEN_2812; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2814 = 10'h2fe == io_inputs_0 ? 7'h0 : _GEN_2813; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2815 = 10'h2ff == io_inputs_0 ? 7'h0 : _GEN_2814; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2816 = 10'h300 == io_inputs_0 ? 7'h0 : _GEN_2815; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2817 = 10'h301 == io_inputs_0 ? 7'h0 : _GEN_2816; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2818 = 10'h302 == io_inputs_0 ? 7'h0 : _GEN_2817; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2819 = 10'h303 == io_inputs_0 ? 7'h0 : _GEN_2818; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2820 = 10'h304 == io_inputs_0 ? 7'h0 : _GEN_2819; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2821 = 10'h305 == io_inputs_0 ? 7'h0 : _GEN_2820; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2822 = 10'h306 == io_inputs_0 ? 7'h0 : _GEN_2821; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2823 = 10'h307 == io_inputs_0 ? 7'h0 : _GEN_2822; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2824 = 10'h308 == io_inputs_0 ? 7'h0 : _GEN_2823; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2825 = 10'h309 == io_inputs_0 ? 7'h0 : _GEN_2824; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2826 = 10'h30a == io_inputs_0 ? 7'h0 : _GEN_2825; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2827 = 10'h30b == io_inputs_0 ? 7'h0 : _GEN_2826; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2828 = 10'h30c == io_inputs_0 ? 7'h0 : _GEN_2827; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2829 = 10'h30d == io_inputs_0 ? 7'h0 : _GEN_2828; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2830 = 10'h30e == io_inputs_0 ? 7'h0 : _GEN_2829; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2831 = 10'h30f == io_inputs_0 ? 7'h0 : _GEN_2830; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2832 = 10'h310 == io_inputs_0 ? 7'h0 : _GEN_2831; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2833 = 10'h311 == io_inputs_0 ? 7'h0 : _GEN_2832; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2834 = 10'h312 == io_inputs_0 ? 7'h0 : _GEN_2833; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2835 = 10'h313 == io_inputs_0 ? 7'h0 : _GEN_2834; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2836 = 10'h314 == io_inputs_0 ? 7'h0 : _GEN_2835; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2837 = 10'h315 == io_inputs_0 ? 7'h0 : _GEN_2836; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2838 = 10'h316 == io_inputs_0 ? 7'h0 : _GEN_2837; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2839 = 10'h317 == io_inputs_0 ? 7'h0 : _GEN_2838; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2840 = 10'h318 == io_inputs_0 ? 7'h0 : _GEN_2839; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2841 = 10'h319 == io_inputs_0 ? 7'h0 : _GEN_2840; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2842 = 10'h31a == io_inputs_0 ? 7'h0 : _GEN_2841; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2843 = 10'h31b == io_inputs_0 ? 7'h0 : _GEN_2842; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2844 = 10'h31c == io_inputs_0 ? 7'h0 : _GEN_2843; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2845 = 10'h31d == io_inputs_0 ? 7'h0 : _GEN_2844; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2846 = 10'h31e == io_inputs_0 ? 7'h0 : _GEN_2845; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2847 = 10'h31f == io_inputs_0 ? 7'h0 : _GEN_2846; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2848 = 10'h320 == io_inputs_0 ? 7'h0 : _GEN_2847; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2849 = 10'h321 == io_inputs_0 ? 7'h0 : _GEN_2848; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2850 = 10'h322 == io_inputs_0 ? 7'h0 : _GEN_2849; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2851 = 10'h323 == io_inputs_0 ? 7'h0 : _GEN_2850; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2852 = 10'h324 == io_inputs_0 ? 7'h0 : _GEN_2851; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2853 = 10'h325 == io_inputs_0 ? 7'h0 : _GEN_2852; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2854 = 10'h326 == io_inputs_0 ? 7'h0 : _GEN_2853; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2855 = 10'h327 == io_inputs_0 ? 7'h0 : _GEN_2854; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2856 = 10'h328 == io_inputs_0 ? 7'h0 : _GEN_2855; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2857 = 10'h329 == io_inputs_0 ? 7'h0 : _GEN_2856; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2858 = 10'h32a == io_inputs_0 ? 7'h0 : _GEN_2857; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2859 = 10'h32b == io_inputs_0 ? 7'h0 : _GEN_2858; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2860 = 10'h32c == io_inputs_0 ? 7'h0 : _GEN_2859; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2861 = 10'h32d == io_inputs_0 ? 7'h0 : _GEN_2860; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2862 = 10'h32e == io_inputs_0 ? 7'h0 : _GEN_2861; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2863 = 10'h32f == io_inputs_0 ? 7'h0 : _GEN_2862; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2864 = 10'h330 == io_inputs_0 ? 7'h0 : _GEN_2863; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2865 = 10'h331 == io_inputs_0 ? 7'h0 : _GEN_2864; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2866 = 10'h332 == io_inputs_0 ? 7'h0 : _GEN_2865; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2867 = 10'h333 == io_inputs_0 ? 7'h0 : _GEN_2866; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2868 = 10'h334 == io_inputs_0 ? 7'h0 : _GEN_2867; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2869 = 10'h335 == io_inputs_0 ? 7'h0 : _GEN_2868; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2870 = 10'h336 == io_inputs_0 ? 7'h0 : _GEN_2869; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2871 = 10'h337 == io_inputs_0 ? 7'h0 : _GEN_2870; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2872 = 10'h338 == io_inputs_0 ? 7'h0 : _GEN_2871; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2873 = 10'h339 == io_inputs_0 ? 7'h0 : _GEN_2872; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2874 = 10'h33a == io_inputs_0 ? 7'h0 : _GEN_2873; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2875 = 10'h33b == io_inputs_0 ? 7'h0 : _GEN_2874; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2876 = 10'h33c == io_inputs_0 ? 7'h0 : _GEN_2875; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2877 = 10'h33d == io_inputs_0 ? 7'h0 : _GEN_2876; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2878 = 10'h33e == io_inputs_0 ? 7'h0 : _GEN_2877; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2879 = 10'h33f == io_inputs_0 ? 7'h0 : _GEN_2878; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2880 = 10'h340 == io_inputs_0 ? 7'h0 : _GEN_2879; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2881 = 10'h341 == io_inputs_0 ? 7'h0 : _GEN_2880; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2882 = 10'h342 == io_inputs_0 ? 7'h0 : _GEN_2881; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2883 = 10'h343 == io_inputs_0 ? 7'h0 : _GEN_2882; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2884 = 10'h344 == io_inputs_0 ? 7'h0 : _GEN_2883; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2885 = 10'h345 == io_inputs_0 ? 7'h0 : _GEN_2884; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2886 = 10'h346 == io_inputs_0 ? 7'h0 : _GEN_2885; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2887 = 10'h347 == io_inputs_0 ? 7'h0 : _GEN_2886; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2888 = 10'h348 == io_inputs_0 ? 7'h0 : _GEN_2887; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2889 = 10'h349 == io_inputs_0 ? 7'h0 : _GEN_2888; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2890 = 10'h34a == io_inputs_0 ? 7'h0 : _GEN_2889; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2891 = 10'h34b == io_inputs_0 ? 7'h0 : _GEN_2890; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2892 = 10'h34c == io_inputs_0 ? 7'h0 : _GEN_2891; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2893 = 10'h34d == io_inputs_0 ? 7'h0 : _GEN_2892; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2894 = 10'h34e == io_inputs_0 ? 7'h0 : _GEN_2893; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2895 = 10'h34f == io_inputs_0 ? 7'h0 : _GEN_2894; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2896 = 10'h350 == io_inputs_0 ? 7'h0 : _GEN_2895; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2897 = 10'h351 == io_inputs_0 ? 7'h0 : _GEN_2896; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2898 = 10'h352 == io_inputs_0 ? 7'h0 : _GEN_2897; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2899 = 10'h353 == io_inputs_0 ? 7'h0 : _GEN_2898; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2900 = 10'h354 == io_inputs_0 ? 7'h0 : _GEN_2899; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2901 = 10'h355 == io_inputs_0 ? 7'h0 : _GEN_2900; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2902 = 10'h356 == io_inputs_0 ? 7'h0 : _GEN_2901; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2903 = 10'h357 == io_inputs_0 ? 7'h0 : _GEN_2902; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2904 = 10'h358 == io_inputs_0 ? 7'h0 : _GEN_2903; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2905 = 10'h359 == io_inputs_0 ? 7'h0 : _GEN_2904; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2906 = 10'h35a == io_inputs_0 ? 7'h0 : _GEN_2905; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2907 = 10'h35b == io_inputs_0 ? 7'h0 : _GEN_2906; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2908 = 10'h35c == io_inputs_0 ? 7'h0 : _GEN_2907; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2909 = 10'h35d == io_inputs_0 ? 7'h0 : _GEN_2908; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2910 = 10'h35e == io_inputs_0 ? 7'h0 : _GEN_2909; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2911 = 10'h35f == io_inputs_0 ? 7'h0 : _GEN_2910; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2912 = 10'h360 == io_inputs_0 ? 7'h0 : _GEN_2911; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2913 = 10'h361 == io_inputs_0 ? 7'h0 : _GEN_2912; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2914 = 10'h362 == io_inputs_0 ? 7'h0 : _GEN_2913; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2915 = 10'h363 == io_inputs_0 ? 7'h0 : _GEN_2914; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2916 = 10'h364 == io_inputs_0 ? 7'h0 : _GEN_2915; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2917 = 10'h365 == io_inputs_0 ? 7'h0 : _GEN_2916; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2918 = 10'h366 == io_inputs_0 ? 7'h0 : _GEN_2917; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2919 = 10'h367 == io_inputs_0 ? 7'h0 : _GEN_2918; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2920 = 10'h368 == io_inputs_0 ? 7'h0 : _GEN_2919; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2921 = 10'h369 == io_inputs_0 ? 7'h0 : _GEN_2920; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2922 = 10'h36a == io_inputs_0 ? 7'h0 : _GEN_2921; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2923 = 10'h36b == io_inputs_0 ? 7'h0 : _GEN_2922; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2924 = 10'h36c == io_inputs_0 ? 7'h0 : _GEN_2923; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2925 = 10'h36d == io_inputs_0 ? 7'h0 : _GEN_2924; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2926 = 10'h36e == io_inputs_0 ? 7'h0 : _GEN_2925; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2927 = 10'h36f == io_inputs_0 ? 7'h0 : _GEN_2926; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2928 = 10'h370 == io_inputs_0 ? 7'h0 : _GEN_2927; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2929 = 10'h371 == io_inputs_0 ? 7'h0 : _GEN_2928; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2930 = 10'h372 == io_inputs_0 ? 7'h0 : _GEN_2929; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2931 = 10'h373 == io_inputs_0 ? 7'h0 : _GEN_2930; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2932 = 10'h374 == io_inputs_0 ? 7'h0 : _GEN_2931; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2933 = 10'h375 == io_inputs_0 ? 7'h0 : _GEN_2932; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2934 = 10'h376 == io_inputs_0 ? 7'h0 : _GEN_2933; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2935 = 10'h377 == io_inputs_0 ? 7'h0 : _GEN_2934; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2936 = 10'h378 == io_inputs_0 ? 7'h0 : _GEN_2935; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2937 = 10'h379 == io_inputs_0 ? 7'h0 : _GEN_2936; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2938 = 10'h37a == io_inputs_0 ? 7'h0 : _GEN_2937; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2939 = 10'h37b == io_inputs_0 ? 7'h0 : _GEN_2938; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2940 = 10'h37c == io_inputs_0 ? 7'h0 : _GEN_2939; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2941 = 10'h37d == io_inputs_0 ? 7'h0 : _GEN_2940; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2942 = 10'h37e == io_inputs_0 ? 7'h0 : _GEN_2941; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2943 = 10'h37f == io_inputs_0 ? 7'h0 : _GEN_2942; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2944 = 10'h380 == io_inputs_0 ? 7'h0 : _GEN_2943; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2945 = 10'h381 == io_inputs_0 ? 7'h0 : _GEN_2944; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2946 = 10'h382 == io_inputs_0 ? 7'h0 : _GEN_2945; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2947 = 10'h383 == io_inputs_0 ? 7'h0 : _GEN_2946; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2948 = 10'h384 == io_inputs_0 ? 7'h0 : _GEN_2947; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2949 = 10'h385 == io_inputs_0 ? 7'h0 : _GEN_2948; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2950 = 10'h386 == io_inputs_0 ? 7'h0 : _GEN_2949; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2951 = 10'h387 == io_inputs_0 ? 7'h0 : _GEN_2950; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2952 = 10'h388 == io_inputs_0 ? 7'h0 : _GEN_2951; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2953 = 10'h389 == io_inputs_0 ? 7'h0 : _GEN_2952; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2954 = 10'h38a == io_inputs_0 ? 7'h0 : _GEN_2953; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2955 = 10'h38b == io_inputs_0 ? 7'h0 : _GEN_2954; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2956 = 10'h38c == io_inputs_0 ? 7'h0 : _GEN_2955; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2957 = 10'h38d == io_inputs_0 ? 7'h0 : _GEN_2956; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2958 = 10'h38e == io_inputs_0 ? 7'h0 : _GEN_2957; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2959 = 10'h38f == io_inputs_0 ? 7'h0 : _GEN_2958; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2960 = 10'h390 == io_inputs_0 ? 7'h0 : _GEN_2959; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2961 = 10'h391 == io_inputs_0 ? 7'h0 : _GEN_2960; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2962 = 10'h392 == io_inputs_0 ? 7'h0 : _GEN_2961; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2963 = 10'h393 == io_inputs_0 ? 7'h0 : _GEN_2962; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2964 = 10'h394 == io_inputs_0 ? 7'h0 : _GEN_2963; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2965 = 10'h395 == io_inputs_0 ? 7'h0 : _GEN_2964; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2966 = 10'h396 == io_inputs_0 ? 7'h0 : _GEN_2965; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2967 = 10'h397 == io_inputs_0 ? 7'h0 : _GEN_2966; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2968 = 10'h398 == io_inputs_0 ? 7'h0 : _GEN_2967; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2969 = 10'h399 == io_inputs_0 ? 7'h0 : _GEN_2968; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2970 = 10'h39a == io_inputs_0 ? 7'h0 : _GEN_2969; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2971 = 10'h39b == io_inputs_0 ? 7'h0 : _GEN_2970; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2972 = 10'h39c == io_inputs_0 ? 7'h0 : _GEN_2971; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2973 = 10'h39d == io_inputs_0 ? 7'h0 : _GEN_2972; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2974 = 10'h39e == io_inputs_0 ? 7'h0 : _GEN_2973; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2975 = 10'h39f == io_inputs_0 ? 7'h0 : _GEN_2974; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2976 = 10'h3a0 == io_inputs_0 ? 7'h0 : _GEN_2975; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2977 = 10'h3a1 == io_inputs_0 ? 7'h0 : _GEN_2976; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2978 = 10'h3a2 == io_inputs_0 ? 7'h0 : _GEN_2977; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2979 = 10'h3a3 == io_inputs_0 ? 7'h0 : _GEN_2978; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2980 = 10'h3a4 == io_inputs_0 ? 7'h0 : _GEN_2979; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2981 = 10'h3a5 == io_inputs_0 ? 7'h0 : _GEN_2980; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2982 = 10'h3a6 == io_inputs_0 ? 7'h0 : _GEN_2981; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2983 = 10'h3a7 == io_inputs_0 ? 7'h0 : _GEN_2982; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2984 = 10'h3a8 == io_inputs_0 ? 7'h0 : _GEN_2983; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2985 = 10'h3a9 == io_inputs_0 ? 7'h0 : _GEN_2984; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2986 = 10'h3aa == io_inputs_0 ? 7'h0 : _GEN_2985; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2987 = 10'h3ab == io_inputs_0 ? 7'h0 : _GEN_2986; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2988 = 10'h3ac == io_inputs_0 ? 7'h0 : _GEN_2987; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2989 = 10'h3ad == io_inputs_0 ? 7'h0 : _GEN_2988; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2990 = 10'h3ae == io_inputs_0 ? 7'h0 : _GEN_2989; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2991 = 10'h3af == io_inputs_0 ? 7'h0 : _GEN_2990; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2992 = 10'h3b0 == io_inputs_0 ? 7'h0 : _GEN_2991; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2993 = 10'h3b1 == io_inputs_0 ? 7'h0 : _GEN_2992; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2994 = 10'h3b2 == io_inputs_0 ? 7'h0 : _GEN_2993; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2995 = 10'h3b3 == io_inputs_0 ? 7'h0 : _GEN_2994; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2996 = 10'h3b4 == io_inputs_0 ? 7'h0 : _GEN_2995; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2997 = 10'h3b5 == io_inputs_0 ? 7'h0 : _GEN_2996; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2998 = 10'h3b6 == io_inputs_0 ? 7'h0 : _GEN_2997; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_2999 = 10'h3b7 == io_inputs_0 ? 7'h0 : _GEN_2998; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3000 = 10'h3b8 == io_inputs_0 ? 7'h0 : _GEN_2999; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3001 = 10'h3b9 == io_inputs_0 ? 7'h0 : _GEN_3000; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3002 = 10'h3ba == io_inputs_0 ? 7'h0 : _GEN_3001; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3003 = 10'h3bb == io_inputs_0 ? 7'h0 : _GEN_3002; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3004 = 10'h3bc == io_inputs_0 ? 7'h0 : _GEN_3003; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3005 = 10'h3bd == io_inputs_0 ? 7'h0 : _GEN_3004; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3006 = 10'h3be == io_inputs_0 ? 7'h0 : _GEN_3005; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3007 = 10'h3bf == io_inputs_0 ? 7'h0 : _GEN_3006; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3008 = 10'h3c0 == io_inputs_0 ? 7'h0 : _GEN_3007; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3009 = 10'h3c1 == io_inputs_0 ? 7'h0 : _GEN_3008; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3010 = 10'h3c2 == io_inputs_0 ? 7'h0 : _GEN_3009; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3011 = 10'h3c3 == io_inputs_0 ? 7'h0 : _GEN_3010; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3012 = 10'h3c4 == io_inputs_0 ? 7'h0 : _GEN_3011; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3013 = 10'h3c5 == io_inputs_0 ? 7'h0 : _GEN_3012; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3014 = 10'h3c6 == io_inputs_0 ? 7'h0 : _GEN_3013; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3015 = 10'h3c7 == io_inputs_0 ? 7'h0 : _GEN_3014; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3016 = 10'h3c8 == io_inputs_0 ? 7'h0 : _GEN_3015; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3017 = 10'h3c9 == io_inputs_0 ? 7'h0 : _GEN_3016; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3018 = 10'h3ca == io_inputs_0 ? 7'h0 : _GEN_3017; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3019 = 10'h3cb == io_inputs_0 ? 7'h0 : _GEN_3018; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3020 = 10'h3cc == io_inputs_0 ? 7'h0 : _GEN_3019; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3021 = 10'h3cd == io_inputs_0 ? 7'h0 : _GEN_3020; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3022 = 10'h3ce == io_inputs_0 ? 7'h0 : _GEN_3021; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3023 = 10'h3cf == io_inputs_0 ? 7'h0 : _GEN_3022; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3024 = 10'h3d0 == io_inputs_0 ? 7'h0 : _GEN_3023; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3025 = 10'h3d1 == io_inputs_0 ? 7'h0 : _GEN_3024; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3026 = 10'h3d2 == io_inputs_0 ? 7'h0 : _GEN_3025; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3027 = 10'h3d3 == io_inputs_0 ? 7'h0 : _GEN_3026; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3028 = 10'h3d4 == io_inputs_0 ? 7'h0 : _GEN_3027; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3029 = 10'h3d5 == io_inputs_0 ? 7'h0 : _GEN_3028; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3030 = 10'h3d6 == io_inputs_0 ? 7'h0 : _GEN_3029; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3031 = 10'h3d7 == io_inputs_0 ? 7'h0 : _GEN_3030; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3032 = 10'h3d8 == io_inputs_0 ? 7'h0 : _GEN_3031; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3033 = 10'h3d9 == io_inputs_0 ? 7'h0 : _GEN_3032; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3034 = 10'h3da == io_inputs_0 ? 7'h0 : _GEN_3033; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3035 = 10'h3db == io_inputs_0 ? 7'h0 : _GEN_3034; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3036 = 10'h3dc == io_inputs_0 ? 7'h0 : _GEN_3035; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3037 = 10'h3dd == io_inputs_0 ? 7'h0 : _GEN_3036; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3038 = 10'h3de == io_inputs_0 ? 7'h0 : _GEN_3037; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3039 = 10'h3df == io_inputs_0 ? 7'h0 : _GEN_3038; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3040 = 10'h3e0 == io_inputs_0 ? 7'h0 : _GEN_3039; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3041 = 10'h3e1 == io_inputs_0 ? 7'h0 : _GEN_3040; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3042 = 10'h3e2 == io_inputs_0 ? 7'h0 : _GEN_3041; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3043 = 10'h3e3 == io_inputs_0 ? 7'h0 : _GEN_3042; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3044 = 10'h3e4 == io_inputs_0 ? 7'h0 : _GEN_3043; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3045 = 10'h3e5 == io_inputs_0 ? 7'h0 : _GEN_3044; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3046 = 10'h3e6 == io_inputs_0 ? 7'h0 : _GEN_3045; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3047 = 10'h3e7 == io_inputs_0 ? 7'h0 : _GEN_3046; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3048 = 10'h3e8 == io_inputs_0 ? 7'h0 : _GEN_3047; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3049 = 10'h3e9 == io_inputs_0 ? 7'h0 : _GEN_3048; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3050 = 10'h3ea == io_inputs_0 ? 7'h0 : _GEN_3049; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3051 = 10'h3eb == io_inputs_0 ? 7'h0 : _GEN_3050; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3052 = 10'h3ec == io_inputs_0 ? 7'h0 : _GEN_3051; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3053 = 10'h3ed == io_inputs_0 ? 7'h0 : _GEN_3052; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3054 = 10'h3ee == io_inputs_0 ? 7'h0 : _GEN_3053; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3055 = 10'h3ef == io_inputs_0 ? 7'h0 : _GEN_3054; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3056 = 10'h3f0 == io_inputs_0 ? 7'h0 : _GEN_3055; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3057 = 10'h3f1 == io_inputs_0 ? 7'h0 : _GEN_3056; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3058 = 10'h3f2 == io_inputs_0 ? 7'h0 : _GEN_3057; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3059 = 10'h3f3 == io_inputs_0 ? 7'h0 : _GEN_3058; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3060 = 10'h3f4 == io_inputs_0 ? 7'h0 : _GEN_3059; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3061 = 10'h3f5 == io_inputs_0 ? 7'h0 : _GEN_3060; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3062 = 10'h3f6 == io_inputs_0 ? 7'h0 : _GEN_3061; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3063 = 10'h3f7 == io_inputs_0 ? 7'h0 : _GEN_3062; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3064 = 10'h3f8 == io_inputs_0 ? 7'h0 : _GEN_3063; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3065 = 10'h3f9 == io_inputs_0 ? 7'h0 : _GEN_3064; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3066 = 10'h3fa == io_inputs_0 ? 7'h0 : _GEN_3065; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3067 = 10'h3fb == io_inputs_0 ? 7'h0 : _GEN_3066; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3068 = 10'h3fc == io_inputs_0 ? 7'h0 : _GEN_3067; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3423 = 10'h15f == io_inputs_0 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3424 = 10'h160 == io_inputs_0 ? 7'h2 : _GEN_3423; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3425 = 10'h161 == io_inputs_0 ? 7'h3 : _GEN_3424; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3426 = 10'h162 == io_inputs_0 ? 7'h4 : _GEN_3425; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3427 = 10'h163 == io_inputs_0 ? 7'h5 : _GEN_3426; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3428 = 10'h164 == io_inputs_0 ? 7'h6 : _GEN_3427; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3429 = 10'h165 == io_inputs_0 ? 7'h7 : _GEN_3428; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3430 = 10'h166 == io_inputs_0 ? 7'h8 : _GEN_3429; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3431 = 10'h167 == io_inputs_0 ? 7'h9 : _GEN_3430; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3432 = 10'h168 == io_inputs_0 ? 7'ha : _GEN_3431; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3433 = 10'h169 == io_inputs_0 ? 7'hb : _GEN_3432; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3434 = 10'h16a == io_inputs_0 ? 7'hc : _GEN_3433; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3435 = 10'h16b == io_inputs_0 ? 7'hd : _GEN_3434; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3436 = 10'h16c == io_inputs_0 ? 7'he : _GEN_3435; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3437 = 10'h16d == io_inputs_0 ? 7'hf : _GEN_3436; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3438 = 10'h16e == io_inputs_0 ? 7'h10 : _GEN_3437; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3439 = 10'h16f == io_inputs_0 ? 7'h11 : _GEN_3438; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3440 = 10'h170 == io_inputs_0 ? 7'h12 : _GEN_3439; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3441 = 10'h171 == io_inputs_0 ? 7'h13 : _GEN_3440; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3442 = 10'h172 == io_inputs_0 ? 7'h14 : _GEN_3441; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3443 = 10'h173 == io_inputs_0 ? 7'h15 : _GEN_3442; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3444 = 10'h174 == io_inputs_0 ? 7'h16 : _GEN_3443; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3445 = 10'h175 == io_inputs_0 ? 7'h17 : _GEN_3444; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3446 = 10'h176 == io_inputs_0 ? 7'h18 : _GEN_3445; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3447 = 10'h177 == io_inputs_0 ? 7'h19 : _GEN_3446; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3448 = 10'h178 == io_inputs_0 ? 7'h1a : _GEN_3447; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3449 = 10'h179 == io_inputs_0 ? 7'h1b : _GEN_3448; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3450 = 10'h17a == io_inputs_0 ? 7'h1c : _GEN_3449; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3451 = 10'h17b == io_inputs_0 ? 7'h1d : _GEN_3450; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3452 = 10'h17c == io_inputs_0 ? 7'h1e : _GEN_3451; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3453 = 10'h17d == io_inputs_0 ? 7'h1f : _GEN_3452; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3454 = 10'h17e == io_inputs_0 ? 7'h20 : _GEN_3453; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3455 = 10'h17f == io_inputs_0 ? 7'h21 : _GEN_3454; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3456 = 10'h180 == io_inputs_0 ? 7'h22 : _GEN_3455; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3457 = 10'h181 == io_inputs_0 ? 7'h23 : _GEN_3456; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3458 = 10'h182 == io_inputs_0 ? 7'h24 : _GEN_3457; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3459 = 10'h183 == io_inputs_0 ? 7'h25 : _GEN_3458; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3460 = 10'h184 == io_inputs_0 ? 7'h26 : _GEN_3459; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3461 = 10'h185 == io_inputs_0 ? 7'h27 : _GEN_3460; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3462 = 10'h186 == io_inputs_0 ? 7'h28 : _GEN_3461; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3463 = 10'h187 == io_inputs_0 ? 7'h29 : _GEN_3462; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3464 = 10'h188 == io_inputs_0 ? 7'h2a : _GEN_3463; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3465 = 10'h189 == io_inputs_0 ? 7'h2b : _GEN_3464; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3466 = 10'h18a == io_inputs_0 ? 7'h2c : _GEN_3465; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3467 = 10'h18b == io_inputs_0 ? 7'h2d : _GEN_3466; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3468 = 10'h18c == io_inputs_0 ? 7'h2e : _GEN_3467; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3469 = 10'h18d == io_inputs_0 ? 7'h2f : _GEN_3468; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3470 = 10'h18e == io_inputs_0 ? 7'h30 : _GEN_3469; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3471 = 10'h18f == io_inputs_0 ? 7'h31 : _GEN_3470; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3472 = 10'h190 == io_inputs_0 ? 7'h32 : _GEN_3471; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3473 = 10'h191 == io_inputs_0 ? 7'h33 : _GEN_3472; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3474 = 10'h192 == io_inputs_0 ? 7'h34 : _GEN_3473; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3475 = 10'h193 == io_inputs_0 ? 7'h35 : _GEN_3474; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3476 = 10'h194 == io_inputs_0 ? 7'h36 : _GEN_3475; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3477 = 10'h195 == io_inputs_0 ? 7'h37 : _GEN_3476; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3478 = 10'h196 == io_inputs_0 ? 7'h38 : _GEN_3477; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3479 = 10'h197 == io_inputs_0 ? 7'h39 : _GEN_3478; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3480 = 10'h198 == io_inputs_0 ? 7'h3a : _GEN_3479; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3481 = 10'h199 == io_inputs_0 ? 7'h3b : _GEN_3480; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3482 = 10'h19a == io_inputs_0 ? 7'h3c : _GEN_3481; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3483 = 10'h19b == io_inputs_0 ? 7'h3d : _GEN_3482; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3484 = 10'h19c == io_inputs_0 ? 7'h3e : _GEN_3483; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3485 = 10'h19d == io_inputs_0 ? 7'h3f : _GEN_3484; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3486 = 10'h19e == io_inputs_0 ? 7'h40 : _GEN_3485; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3487 = 10'h19f == io_inputs_0 ? 7'h41 : _GEN_3486; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3488 = 10'h1a0 == io_inputs_0 ? 7'h42 : _GEN_3487; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3489 = 10'h1a1 == io_inputs_0 ? 7'h43 : _GEN_3488; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3490 = 10'h1a2 == io_inputs_0 ? 7'h44 : _GEN_3489; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3491 = 10'h1a3 == io_inputs_0 ? 7'h45 : _GEN_3490; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3492 = 10'h1a4 == io_inputs_0 ? 7'h46 : _GEN_3491; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3493 = 10'h1a5 == io_inputs_0 ? 7'h47 : _GEN_3492; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3494 = 10'h1a6 == io_inputs_0 ? 7'h48 : _GEN_3493; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3495 = 10'h1a7 == io_inputs_0 ? 7'h49 : _GEN_3494; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3496 = 10'h1a8 == io_inputs_0 ? 7'h4a : _GEN_3495; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3497 = 10'h1a9 == io_inputs_0 ? 7'h4b : _GEN_3496; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3498 = 10'h1aa == io_inputs_0 ? 7'h4c : _GEN_3497; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3499 = 10'h1ab == io_inputs_0 ? 7'h4d : _GEN_3498; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3500 = 10'h1ac == io_inputs_0 ? 7'h4e : _GEN_3499; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3501 = 10'h1ad == io_inputs_0 ? 7'h4f : _GEN_3500; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3502 = 10'h1ae == io_inputs_0 ? 7'h50 : _GEN_3501; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3503 = 10'h1af == io_inputs_0 ? 7'h51 : _GEN_3502; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3504 = 10'h1b0 == io_inputs_0 ? 7'h52 : _GEN_3503; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3505 = 10'h1b1 == io_inputs_0 ? 7'h53 : _GEN_3504; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3506 = 10'h1b2 == io_inputs_0 ? 7'h54 : _GEN_3505; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3507 = 10'h1b3 == io_inputs_0 ? 7'h55 : _GEN_3506; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3508 = 10'h1b4 == io_inputs_0 ? 7'h56 : _GEN_3507; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3509 = 10'h1b5 == io_inputs_0 ? 7'h57 : _GEN_3508; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3510 = 10'h1b6 == io_inputs_0 ? 7'h58 : _GEN_3509; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3511 = 10'h1b7 == io_inputs_0 ? 7'h59 : _GEN_3510; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3512 = 10'h1b8 == io_inputs_0 ? 7'h5a : _GEN_3511; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3513 = 10'h1b9 == io_inputs_0 ? 7'h5b : _GEN_3512; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3514 = 10'h1ba == io_inputs_0 ? 7'h5c : _GEN_3513; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3515 = 10'h1bb == io_inputs_0 ? 7'h5d : _GEN_3514; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3516 = 10'h1bc == io_inputs_0 ? 7'h5e : _GEN_3515; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3517 = 10'h1bd == io_inputs_0 ? 7'h5f : _GEN_3516; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3518 = 10'h1be == io_inputs_0 ? 7'h60 : _GEN_3517; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3519 = 10'h1bf == io_inputs_0 ? 7'h61 : _GEN_3518; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3520 = 10'h1c0 == io_inputs_0 ? 7'h62 : _GEN_3519; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3521 = 10'h1c1 == io_inputs_0 ? 7'h63 : _GEN_3520; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3522 = 10'h1c2 == io_inputs_0 ? 7'h64 : _GEN_3521; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3523 = 10'h1c3 == io_inputs_0 ? 7'h63 : _GEN_3522; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3524 = 10'h1c4 == io_inputs_0 ? 7'h62 : _GEN_3523; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3525 = 10'h1c5 == io_inputs_0 ? 7'h61 : _GEN_3524; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3526 = 10'h1c6 == io_inputs_0 ? 7'h60 : _GEN_3525; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3527 = 10'h1c7 == io_inputs_0 ? 7'h5f : _GEN_3526; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3528 = 10'h1c8 == io_inputs_0 ? 7'h5e : _GEN_3527; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3529 = 10'h1c9 == io_inputs_0 ? 7'h5d : _GEN_3528; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3530 = 10'h1ca == io_inputs_0 ? 7'h5c : _GEN_3529; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3531 = 10'h1cb == io_inputs_0 ? 7'h5b : _GEN_3530; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3532 = 10'h1cc == io_inputs_0 ? 7'h5a : _GEN_3531; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3533 = 10'h1cd == io_inputs_0 ? 7'h59 : _GEN_3532; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3534 = 10'h1ce == io_inputs_0 ? 7'h58 : _GEN_3533; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3535 = 10'h1cf == io_inputs_0 ? 7'h57 : _GEN_3534; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3536 = 10'h1d0 == io_inputs_0 ? 7'h56 : _GEN_3535; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3537 = 10'h1d1 == io_inputs_0 ? 7'h55 : _GEN_3536; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3538 = 10'h1d2 == io_inputs_0 ? 7'h54 : _GEN_3537; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3539 = 10'h1d3 == io_inputs_0 ? 7'h53 : _GEN_3538; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3540 = 10'h1d4 == io_inputs_0 ? 7'h52 : _GEN_3539; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3541 = 10'h1d5 == io_inputs_0 ? 7'h51 : _GEN_3540; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3542 = 10'h1d6 == io_inputs_0 ? 7'h50 : _GEN_3541; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3543 = 10'h1d7 == io_inputs_0 ? 7'h4f : _GEN_3542; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3544 = 10'h1d8 == io_inputs_0 ? 7'h4e : _GEN_3543; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3545 = 10'h1d9 == io_inputs_0 ? 7'h4d : _GEN_3544; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3546 = 10'h1da == io_inputs_0 ? 7'h4c : _GEN_3545; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3547 = 10'h1db == io_inputs_0 ? 7'h4b : _GEN_3546; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3548 = 10'h1dc == io_inputs_0 ? 7'h4a : _GEN_3547; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3549 = 10'h1dd == io_inputs_0 ? 7'h49 : _GEN_3548; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3550 = 10'h1de == io_inputs_0 ? 7'h48 : _GEN_3549; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3551 = 10'h1df == io_inputs_0 ? 7'h47 : _GEN_3550; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3552 = 10'h1e0 == io_inputs_0 ? 7'h46 : _GEN_3551; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3553 = 10'h1e1 == io_inputs_0 ? 7'h45 : _GEN_3552; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3554 = 10'h1e2 == io_inputs_0 ? 7'h44 : _GEN_3553; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3555 = 10'h1e3 == io_inputs_0 ? 7'h43 : _GEN_3554; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3556 = 10'h1e4 == io_inputs_0 ? 7'h42 : _GEN_3555; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3557 = 10'h1e5 == io_inputs_0 ? 7'h41 : _GEN_3556; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3558 = 10'h1e6 == io_inputs_0 ? 7'h40 : _GEN_3557; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3559 = 10'h1e7 == io_inputs_0 ? 7'h3f : _GEN_3558; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3560 = 10'h1e8 == io_inputs_0 ? 7'h3e : _GEN_3559; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3561 = 10'h1e9 == io_inputs_0 ? 7'h3d : _GEN_3560; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3562 = 10'h1ea == io_inputs_0 ? 7'h3c : _GEN_3561; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3563 = 10'h1eb == io_inputs_0 ? 7'h3b : _GEN_3562; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3564 = 10'h1ec == io_inputs_0 ? 7'h3a : _GEN_3563; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3565 = 10'h1ed == io_inputs_0 ? 7'h39 : _GEN_3564; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3566 = 10'h1ee == io_inputs_0 ? 7'h38 : _GEN_3565; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3567 = 10'h1ef == io_inputs_0 ? 7'h37 : _GEN_3566; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3568 = 10'h1f0 == io_inputs_0 ? 7'h36 : _GEN_3567; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3569 = 10'h1f1 == io_inputs_0 ? 7'h35 : _GEN_3568; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3570 = 10'h1f2 == io_inputs_0 ? 7'h34 : _GEN_3569; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3571 = 10'h1f3 == io_inputs_0 ? 7'h33 : _GEN_3570; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3572 = 10'h1f4 == io_inputs_0 ? 7'h32 : _GEN_3571; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3573 = 10'h1f5 == io_inputs_0 ? 7'h31 : _GEN_3572; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3574 = 10'h1f6 == io_inputs_0 ? 7'h30 : _GEN_3573; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3575 = 10'h1f7 == io_inputs_0 ? 7'h2f : _GEN_3574; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3576 = 10'h1f8 == io_inputs_0 ? 7'h2e : _GEN_3575; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3577 = 10'h1f9 == io_inputs_0 ? 7'h2d : _GEN_3576; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3578 = 10'h1fa == io_inputs_0 ? 7'h2c : _GEN_3577; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3579 = 10'h1fb == io_inputs_0 ? 7'h2b : _GEN_3578; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3580 = 10'h1fc == io_inputs_0 ? 7'h2a : _GEN_3579; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3581 = 10'h1fd == io_inputs_0 ? 7'h29 : _GEN_3580; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3582 = 10'h1fe == io_inputs_0 ? 7'h28 : _GEN_3581; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3583 = 10'h1ff == io_inputs_0 ? 7'h27 : _GEN_3582; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3584 = 10'h200 == io_inputs_0 ? 7'h26 : _GEN_3583; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3585 = 10'h201 == io_inputs_0 ? 7'h25 : _GEN_3584; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3586 = 10'h202 == io_inputs_0 ? 7'h24 : _GEN_3585; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3587 = 10'h203 == io_inputs_0 ? 7'h23 : _GEN_3586; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3588 = 10'h204 == io_inputs_0 ? 7'h22 : _GEN_3587; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3589 = 10'h205 == io_inputs_0 ? 7'h21 : _GEN_3588; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3590 = 10'h206 == io_inputs_0 ? 7'h20 : _GEN_3589; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3591 = 10'h207 == io_inputs_0 ? 7'h1f : _GEN_3590; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3592 = 10'h208 == io_inputs_0 ? 7'h1e : _GEN_3591; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3593 = 10'h209 == io_inputs_0 ? 7'h1d : _GEN_3592; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3594 = 10'h20a == io_inputs_0 ? 7'h1c : _GEN_3593; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3595 = 10'h20b == io_inputs_0 ? 7'h1b : _GEN_3594; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3596 = 10'h20c == io_inputs_0 ? 7'h1a : _GEN_3595; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3597 = 10'h20d == io_inputs_0 ? 7'h19 : _GEN_3596; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3598 = 10'h20e == io_inputs_0 ? 7'h18 : _GEN_3597; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3599 = 10'h20f == io_inputs_0 ? 7'h17 : _GEN_3598; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3600 = 10'h210 == io_inputs_0 ? 7'h16 : _GEN_3599; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3601 = 10'h211 == io_inputs_0 ? 7'h15 : _GEN_3600; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3602 = 10'h212 == io_inputs_0 ? 7'h14 : _GEN_3601; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3603 = 10'h213 == io_inputs_0 ? 7'h13 : _GEN_3602; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3604 = 10'h214 == io_inputs_0 ? 7'h12 : _GEN_3603; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3605 = 10'h215 == io_inputs_0 ? 7'h11 : _GEN_3604; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3606 = 10'h216 == io_inputs_0 ? 7'h10 : _GEN_3605; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3607 = 10'h217 == io_inputs_0 ? 7'hf : _GEN_3606; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3608 = 10'h218 == io_inputs_0 ? 7'he : _GEN_3607; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3609 = 10'h219 == io_inputs_0 ? 7'hd : _GEN_3608; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3610 = 10'h21a == io_inputs_0 ? 7'hc : _GEN_3609; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3611 = 10'h21b == io_inputs_0 ? 7'hb : _GEN_3610; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3612 = 10'h21c == io_inputs_0 ? 7'ha : _GEN_3611; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3613 = 10'h21d == io_inputs_0 ? 7'h9 : _GEN_3612; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3614 = 10'h21e == io_inputs_0 ? 7'h8 : _GEN_3613; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3615 = 10'h21f == io_inputs_0 ? 7'h7 : _GEN_3614; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3616 = 10'h220 == io_inputs_0 ? 7'h6 : _GEN_3615; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3617 = 10'h221 == io_inputs_0 ? 7'h5 : _GEN_3616; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3618 = 10'h222 == io_inputs_0 ? 7'h4 : _GEN_3617; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3619 = 10'h223 == io_inputs_0 ? 7'h3 : _GEN_3618; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3620 = 10'h224 == io_inputs_0 ? 7'h2 : _GEN_3619; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3621 = 10'h225 == io_inputs_0 ? 7'h1 : _GEN_3620; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3622 = 10'h226 == io_inputs_0 ? 7'h0 : _GEN_3621; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3623 = 10'h227 == io_inputs_0 ? 7'h0 : _GEN_3622; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3624 = 10'h228 == io_inputs_0 ? 7'h0 : _GEN_3623; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3625 = 10'h229 == io_inputs_0 ? 7'h0 : _GEN_3624; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3626 = 10'h22a == io_inputs_0 ? 7'h0 : _GEN_3625; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3627 = 10'h22b == io_inputs_0 ? 7'h0 : _GEN_3626; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3628 = 10'h22c == io_inputs_0 ? 7'h0 : _GEN_3627; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3629 = 10'h22d == io_inputs_0 ? 7'h0 : _GEN_3628; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3630 = 10'h22e == io_inputs_0 ? 7'h0 : _GEN_3629; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3631 = 10'h22f == io_inputs_0 ? 7'h0 : _GEN_3630; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3632 = 10'h230 == io_inputs_0 ? 7'h0 : _GEN_3631; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3633 = 10'h231 == io_inputs_0 ? 7'h0 : _GEN_3632; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3634 = 10'h232 == io_inputs_0 ? 7'h0 : _GEN_3633; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3635 = 10'h233 == io_inputs_0 ? 7'h0 : _GEN_3634; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3636 = 10'h234 == io_inputs_0 ? 7'h0 : _GEN_3635; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3637 = 10'h235 == io_inputs_0 ? 7'h0 : _GEN_3636; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3638 = 10'h236 == io_inputs_0 ? 7'h0 : _GEN_3637; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3639 = 10'h237 == io_inputs_0 ? 7'h0 : _GEN_3638; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3640 = 10'h238 == io_inputs_0 ? 7'h0 : _GEN_3639; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3641 = 10'h239 == io_inputs_0 ? 7'h0 : _GEN_3640; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3642 = 10'h23a == io_inputs_0 ? 7'h0 : _GEN_3641; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3643 = 10'h23b == io_inputs_0 ? 7'h0 : _GEN_3642; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3644 = 10'h23c == io_inputs_0 ? 7'h0 : _GEN_3643; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3645 = 10'h23d == io_inputs_0 ? 7'h0 : _GEN_3644; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3646 = 10'h23e == io_inputs_0 ? 7'h0 : _GEN_3645; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3647 = 10'h23f == io_inputs_0 ? 7'h0 : _GEN_3646; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3648 = 10'h240 == io_inputs_0 ? 7'h0 : _GEN_3647; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3649 = 10'h241 == io_inputs_0 ? 7'h0 : _GEN_3648; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3650 = 10'h242 == io_inputs_0 ? 7'h0 : _GEN_3649; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3651 = 10'h243 == io_inputs_0 ? 7'h0 : _GEN_3650; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3652 = 10'h244 == io_inputs_0 ? 7'h0 : _GEN_3651; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3653 = 10'h245 == io_inputs_0 ? 7'h0 : _GEN_3652; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3654 = 10'h246 == io_inputs_0 ? 7'h0 : _GEN_3653; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3655 = 10'h247 == io_inputs_0 ? 7'h0 : _GEN_3654; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3656 = 10'h248 == io_inputs_0 ? 7'h0 : _GEN_3655; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3657 = 10'h249 == io_inputs_0 ? 7'h0 : _GEN_3656; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3658 = 10'h24a == io_inputs_0 ? 7'h0 : _GEN_3657; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3659 = 10'h24b == io_inputs_0 ? 7'h0 : _GEN_3658; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3660 = 10'h24c == io_inputs_0 ? 7'h0 : _GEN_3659; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3661 = 10'h24d == io_inputs_0 ? 7'h0 : _GEN_3660; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3662 = 10'h24e == io_inputs_0 ? 7'h0 : _GEN_3661; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3663 = 10'h24f == io_inputs_0 ? 7'h0 : _GEN_3662; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3664 = 10'h250 == io_inputs_0 ? 7'h0 : _GEN_3663; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3665 = 10'h251 == io_inputs_0 ? 7'h0 : _GEN_3664; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3666 = 10'h252 == io_inputs_0 ? 7'h0 : _GEN_3665; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3667 = 10'h253 == io_inputs_0 ? 7'h0 : _GEN_3666; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3668 = 10'h254 == io_inputs_0 ? 7'h0 : _GEN_3667; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3669 = 10'h255 == io_inputs_0 ? 7'h0 : _GEN_3668; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3670 = 10'h256 == io_inputs_0 ? 7'h0 : _GEN_3669; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3671 = 10'h257 == io_inputs_0 ? 7'h0 : _GEN_3670; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3672 = 10'h258 == io_inputs_0 ? 7'h0 : _GEN_3671; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3673 = 10'h259 == io_inputs_0 ? 7'h0 : _GEN_3672; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3674 = 10'h25a == io_inputs_0 ? 7'h0 : _GEN_3673; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3675 = 10'h25b == io_inputs_0 ? 7'h0 : _GEN_3674; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3676 = 10'h25c == io_inputs_0 ? 7'h0 : _GEN_3675; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3677 = 10'h25d == io_inputs_0 ? 7'h0 : _GEN_3676; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3678 = 10'h25e == io_inputs_0 ? 7'h0 : _GEN_3677; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3679 = 10'h25f == io_inputs_0 ? 7'h0 : _GEN_3678; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3680 = 10'h260 == io_inputs_0 ? 7'h0 : _GEN_3679; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3681 = 10'h261 == io_inputs_0 ? 7'h0 : _GEN_3680; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3682 = 10'h262 == io_inputs_0 ? 7'h0 : _GEN_3681; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3683 = 10'h263 == io_inputs_0 ? 7'h0 : _GEN_3682; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3684 = 10'h264 == io_inputs_0 ? 7'h0 : _GEN_3683; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3685 = 10'h265 == io_inputs_0 ? 7'h0 : _GEN_3684; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3686 = 10'h266 == io_inputs_0 ? 7'h0 : _GEN_3685; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3687 = 10'h267 == io_inputs_0 ? 7'h0 : _GEN_3686; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3688 = 10'h268 == io_inputs_0 ? 7'h0 : _GEN_3687; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3689 = 10'h269 == io_inputs_0 ? 7'h0 : _GEN_3688; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3690 = 10'h26a == io_inputs_0 ? 7'h0 : _GEN_3689; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3691 = 10'h26b == io_inputs_0 ? 7'h0 : _GEN_3690; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3692 = 10'h26c == io_inputs_0 ? 7'h0 : _GEN_3691; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3693 = 10'h26d == io_inputs_0 ? 7'h0 : _GEN_3692; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3694 = 10'h26e == io_inputs_0 ? 7'h0 : _GEN_3693; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3695 = 10'h26f == io_inputs_0 ? 7'h0 : _GEN_3694; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3696 = 10'h270 == io_inputs_0 ? 7'h0 : _GEN_3695; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3697 = 10'h271 == io_inputs_0 ? 7'h0 : _GEN_3696; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3698 = 10'h272 == io_inputs_0 ? 7'h0 : _GEN_3697; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3699 = 10'h273 == io_inputs_0 ? 7'h0 : _GEN_3698; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3700 = 10'h274 == io_inputs_0 ? 7'h0 : _GEN_3699; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3701 = 10'h275 == io_inputs_0 ? 7'h0 : _GEN_3700; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3702 = 10'h276 == io_inputs_0 ? 7'h0 : _GEN_3701; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3703 = 10'h277 == io_inputs_0 ? 7'h0 : _GEN_3702; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3704 = 10'h278 == io_inputs_0 ? 7'h0 : _GEN_3703; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3705 = 10'h279 == io_inputs_0 ? 7'h0 : _GEN_3704; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3706 = 10'h27a == io_inputs_0 ? 7'h0 : _GEN_3705; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3707 = 10'h27b == io_inputs_0 ? 7'h0 : _GEN_3706; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3708 = 10'h27c == io_inputs_0 ? 7'h0 : _GEN_3707; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3709 = 10'h27d == io_inputs_0 ? 7'h0 : _GEN_3708; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3710 = 10'h27e == io_inputs_0 ? 7'h0 : _GEN_3709; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3711 = 10'h27f == io_inputs_0 ? 7'h0 : _GEN_3710; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3712 = 10'h280 == io_inputs_0 ? 7'h0 : _GEN_3711; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3713 = 10'h281 == io_inputs_0 ? 7'h0 : _GEN_3712; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3714 = 10'h282 == io_inputs_0 ? 7'h0 : _GEN_3713; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3715 = 10'h283 == io_inputs_0 ? 7'h0 : _GEN_3714; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3716 = 10'h284 == io_inputs_0 ? 7'h0 : _GEN_3715; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3717 = 10'h285 == io_inputs_0 ? 7'h0 : _GEN_3716; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3718 = 10'h286 == io_inputs_0 ? 7'h0 : _GEN_3717; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3719 = 10'h287 == io_inputs_0 ? 7'h0 : _GEN_3718; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3720 = 10'h288 == io_inputs_0 ? 7'h0 : _GEN_3719; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3721 = 10'h289 == io_inputs_0 ? 7'h0 : _GEN_3720; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3722 = 10'h28a == io_inputs_0 ? 7'h0 : _GEN_3721; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3723 = 10'h28b == io_inputs_0 ? 7'h0 : _GEN_3722; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3724 = 10'h28c == io_inputs_0 ? 7'h0 : _GEN_3723; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3725 = 10'h28d == io_inputs_0 ? 7'h0 : _GEN_3724; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3726 = 10'h28e == io_inputs_0 ? 7'h0 : _GEN_3725; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3727 = 10'h28f == io_inputs_0 ? 7'h0 : _GEN_3726; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3728 = 10'h290 == io_inputs_0 ? 7'h0 : _GEN_3727; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3729 = 10'h291 == io_inputs_0 ? 7'h0 : _GEN_3728; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3730 = 10'h292 == io_inputs_0 ? 7'h0 : _GEN_3729; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3731 = 10'h293 == io_inputs_0 ? 7'h0 : _GEN_3730; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3732 = 10'h294 == io_inputs_0 ? 7'h0 : _GEN_3731; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3733 = 10'h295 == io_inputs_0 ? 7'h0 : _GEN_3732; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3734 = 10'h296 == io_inputs_0 ? 7'h0 : _GEN_3733; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3735 = 10'h297 == io_inputs_0 ? 7'h0 : _GEN_3734; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3736 = 10'h298 == io_inputs_0 ? 7'h0 : _GEN_3735; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3737 = 10'h299 == io_inputs_0 ? 7'h0 : _GEN_3736; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3738 = 10'h29a == io_inputs_0 ? 7'h0 : _GEN_3737; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3739 = 10'h29b == io_inputs_0 ? 7'h0 : _GEN_3738; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3740 = 10'h29c == io_inputs_0 ? 7'h0 : _GEN_3739; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3741 = 10'h29d == io_inputs_0 ? 7'h0 : _GEN_3740; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3742 = 10'h29e == io_inputs_0 ? 7'h0 : _GEN_3741; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3743 = 10'h29f == io_inputs_0 ? 7'h0 : _GEN_3742; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3744 = 10'h2a0 == io_inputs_0 ? 7'h0 : _GEN_3743; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3745 = 10'h2a1 == io_inputs_0 ? 7'h0 : _GEN_3744; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3746 = 10'h2a2 == io_inputs_0 ? 7'h0 : _GEN_3745; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3747 = 10'h2a3 == io_inputs_0 ? 7'h0 : _GEN_3746; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3748 = 10'h2a4 == io_inputs_0 ? 7'h0 : _GEN_3747; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3749 = 10'h2a5 == io_inputs_0 ? 7'h0 : _GEN_3748; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3750 = 10'h2a6 == io_inputs_0 ? 7'h0 : _GEN_3749; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3751 = 10'h2a7 == io_inputs_0 ? 7'h0 : _GEN_3750; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3752 = 10'h2a8 == io_inputs_0 ? 7'h0 : _GEN_3751; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3753 = 10'h2a9 == io_inputs_0 ? 7'h0 : _GEN_3752; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3754 = 10'h2aa == io_inputs_0 ? 7'h0 : _GEN_3753; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3755 = 10'h2ab == io_inputs_0 ? 7'h0 : _GEN_3754; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3756 = 10'h2ac == io_inputs_0 ? 7'h0 : _GEN_3755; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3757 = 10'h2ad == io_inputs_0 ? 7'h0 : _GEN_3756; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3758 = 10'h2ae == io_inputs_0 ? 7'h0 : _GEN_3757; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3759 = 10'h2af == io_inputs_0 ? 7'h0 : _GEN_3758; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3760 = 10'h2b0 == io_inputs_0 ? 7'h0 : _GEN_3759; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3761 = 10'h2b1 == io_inputs_0 ? 7'h0 : _GEN_3760; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3762 = 10'h2b2 == io_inputs_0 ? 7'h0 : _GEN_3761; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3763 = 10'h2b3 == io_inputs_0 ? 7'h0 : _GEN_3762; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3764 = 10'h2b4 == io_inputs_0 ? 7'h0 : _GEN_3763; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3765 = 10'h2b5 == io_inputs_0 ? 7'h0 : _GEN_3764; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3766 = 10'h2b6 == io_inputs_0 ? 7'h0 : _GEN_3765; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3767 = 10'h2b7 == io_inputs_0 ? 7'h0 : _GEN_3766; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3768 = 10'h2b8 == io_inputs_0 ? 7'h0 : _GEN_3767; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3769 = 10'h2b9 == io_inputs_0 ? 7'h0 : _GEN_3768; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3770 = 10'h2ba == io_inputs_0 ? 7'h0 : _GEN_3769; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3771 = 10'h2bb == io_inputs_0 ? 7'h0 : _GEN_3770; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3772 = 10'h2bc == io_inputs_0 ? 7'h0 : _GEN_3771; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3773 = 10'h2bd == io_inputs_0 ? 7'h0 : _GEN_3772; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3774 = 10'h2be == io_inputs_0 ? 7'h0 : _GEN_3773; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3775 = 10'h2bf == io_inputs_0 ? 7'h0 : _GEN_3774; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3776 = 10'h2c0 == io_inputs_0 ? 7'h0 : _GEN_3775; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3777 = 10'h2c1 == io_inputs_0 ? 7'h0 : _GEN_3776; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3778 = 10'h2c2 == io_inputs_0 ? 7'h0 : _GEN_3777; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3779 = 10'h2c3 == io_inputs_0 ? 7'h0 : _GEN_3778; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3780 = 10'h2c4 == io_inputs_0 ? 7'h0 : _GEN_3779; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3781 = 10'h2c5 == io_inputs_0 ? 7'h0 : _GEN_3780; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3782 = 10'h2c6 == io_inputs_0 ? 7'h0 : _GEN_3781; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3783 = 10'h2c7 == io_inputs_0 ? 7'h0 : _GEN_3782; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3784 = 10'h2c8 == io_inputs_0 ? 7'h0 : _GEN_3783; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3785 = 10'h2c9 == io_inputs_0 ? 7'h0 : _GEN_3784; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3786 = 10'h2ca == io_inputs_0 ? 7'h0 : _GEN_3785; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3787 = 10'h2cb == io_inputs_0 ? 7'h0 : _GEN_3786; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3788 = 10'h2cc == io_inputs_0 ? 7'h0 : _GEN_3787; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3789 = 10'h2cd == io_inputs_0 ? 7'h0 : _GEN_3788; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3790 = 10'h2ce == io_inputs_0 ? 7'h0 : _GEN_3789; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3791 = 10'h2cf == io_inputs_0 ? 7'h0 : _GEN_3790; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3792 = 10'h2d0 == io_inputs_0 ? 7'h0 : _GEN_3791; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3793 = 10'h2d1 == io_inputs_0 ? 7'h0 : _GEN_3792; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3794 = 10'h2d2 == io_inputs_0 ? 7'h0 : _GEN_3793; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3795 = 10'h2d3 == io_inputs_0 ? 7'h0 : _GEN_3794; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3796 = 10'h2d4 == io_inputs_0 ? 7'h0 : _GEN_3795; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3797 = 10'h2d5 == io_inputs_0 ? 7'h0 : _GEN_3796; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3798 = 10'h2d6 == io_inputs_0 ? 7'h0 : _GEN_3797; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3799 = 10'h2d7 == io_inputs_0 ? 7'h0 : _GEN_3798; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3800 = 10'h2d8 == io_inputs_0 ? 7'h0 : _GEN_3799; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3801 = 10'h2d9 == io_inputs_0 ? 7'h0 : _GEN_3800; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3802 = 10'h2da == io_inputs_0 ? 7'h0 : _GEN_3801; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3803 = 10'h2db == io_inputs_0 ? 7'h0 : _GEN_3802; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3804 = 10'h2dc == io_inputs_0 ? 7'h0 : _GEN_3803; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3805 = 10'h2dd == io_inputs_0 ? 7'h0 : _GEN_3804; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3806 = 10'h2de == io_inputs_0 ? 7'h0 : _GEN_3805; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3807 = 10'h2df == io_inputs_0 ? 7'h0 : _GEN_3806; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3808 = 10'h2e0 == io_inputs_0 ? 7'h0 : _GEN_3807; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3809 = 10'h2e1 == io_inputs_0 ? 7'h0 : _GEN_3808; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3810 = 10'h2e2 == io_inputs_0 ? 7'h0 : _GEN_3809; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3811 = 10'h2e3 == io_inputs_0 ? 7'h0 : _GEN_3810; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3812 = 10'h2e4 == io_inputs_0 ? 7'h0 : _GEN_3811; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3813 = 10'h2e5 == io_inputs_0 ? 7'h0 : _GEN_3812; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3814 = 10'h2e6 == io_inputs_0 ? 7'h0 : _GEN_3813; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3815 = 10'h2e7 == io_inputs_0 ? 7'h0 : _GEN_3814; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3816 = 10'h2e8 == io_inputs_0 ? 7'h0 : _GEN_3815; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3817 = 10'h2e9 == io_inputs_0 ? 7'h0 : _GEN_3816; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3818 = 10'h2ea == io_inputs_0 ? 7'h0 : _GEN_3817; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3819 = 10'h2eb == io_inputs_0 ? 7'h0 : _GEN_3818; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3820 = 10'h2ec == io_inputs_0 ? 7'h0 : _GEN_3819; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3821 = 10'h2ed == io_inputs_0 ? 7'h0 : _GEN_3820; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3822 = 10'h2ee == io_inputs_0 ? 7'h0 : _GEN_3821; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3823 = 10'h2ef == io_inputs_0 ? 7'h0 : _GEN_3822; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3824 = 10'h2f0 == io_inputs_0 ? 7'h0 : _GEN_3823; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3825 = 10'h2f1 == io_inputs_0 ? 7'h0 : _GEN_3824; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3826 = 10'h2f2 == io_inputs_0 ? 7'h0 : _GEN_3825; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3827 = 10'h2f3 == io_inputs_0 ? 7'h0 : _GEN_3826; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3828 = 10'h2f4 == io_inputs_0 ? 7'h0 : _GEN_3827; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3829 = 10'h2f5 == io_inputs_0 ? 7'h0 : _GEN_3828; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3830 = 10'h2f6 == io_inputs_0 ? 7'h0 : _GEN_3829; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3831 = 10'h2f7 == io_inputs_0 ? 7'h0 : _GEN_3830; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3832 = 10'h2f8 == io_inputs_0 ? 7'h0 : _GEN_3831; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3833 = 10'h2f9 == io_inputs_0 ? 7'h0 : _GEN_3832; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3834 = 10'h2fa == io_inputs_0 ? 7'h0 : _GEN_3833; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3835 = 10'h2fb == io_inputs_0 ? 7'h0 : _GEN_3834; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3836 = 10'h2fc == io_inputs_0 ? 7'h0 : _GEN_3835; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3837 = 10'h2fd == io_inputs_0 ? 7'h0 : _GEN_3836; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3838 = 10'h2fe == io_inputs_0 ? 7'h0 : _GEN_3837; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3839 = 10'h2ff == io_inputs_0 ? 7'h0 : _GEN_3838; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3840 = 10'h300 == io_inputs_0 ? 7'h0 : _GEN_3839; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3841 = 10'h301 == io_inputs_0 ? 7'h0 : _GEN_3840; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3842 = 10'h302 == io_inputs_0 ? 7'h0 : _GEN_3841; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3843 = 10'h303 == io_inputs_0 ? 7'h0 : _GEN_3842; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3844 = 10'h304 == io_inputs_0 ? 7'h0 : _GEN_3843; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3845 = 10'h305 == io_inputs_0 ? 7'h0 : _GEN_3844; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3846 = 10'h306 == io_inputs_0 ? 7'h0 : _GEN_3845; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3847 = 10'h307 == io_inputs_0 ? 7'h0 : _GEN_3846; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3848 = 10'h308 == io_inputs_0 ? 7'h0 : _GEN_3847; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3849 = 10'h309 == io_inputs_0 ? 7'h0 : _GEN_3848; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3850 = 10'h30a == io_inputs_0 ? 7'h0 : _GEN_3849; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3851 = 10'h30b == io_inputs_0 ? 7'h0 : _GEN_3850; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3852 = 10'h30c == io_inputs_0 ? 7'h0 : _GEN_3851; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3853 = 10'h30d == io_inputs_0 ? 7'h0 : _GEN_3852; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3854 = 10'h30e == io_inputs_0 ? 7'h0 : _GEN_3853; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3855 = 10'h30f == io_inputs_0 ? 7'h0 : _GEN_3854; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3856 = 10'h310 == io_inputs_0 ? 7'h0 : _GEN_3855; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3857 = 10'h311 == io_inputs_0 ? 7'h0 : _GEN_3856; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3858 = 10'h312 == io_inputs_0 ? 7'h0 : _GEN_3857; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3859 = 10'h313 == io_inputs_0 ? 7'h0 : _GEN_3858; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3860 = 10'h314 == io_inputs_0 ? 7'h0 : _GEN_3859; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3861 = 10'h315 == io_inputs_0 ? 7'h0 : _GEN_3860; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3862 = 10'h316 == io_inputs_0 ? 7'h0 : _GEN_3861; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3863 = 10'h317 == io_inputs_0 ? 7'h0 : _GEN_3862; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3864 = 10'h318 == io_inputs_0 ? 7'h0 : _GEN_3863; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3865 = 10'h319 == io_inputs_0 ? 7'h0 : _GEN_3864; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3866 = 10'h31a == io_inputs_0 ? 7'h0 : _GEN_3865; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3867 = 10'h31b == io_inputs_0 ? 7'h0 : _GEN_3866; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3868 = 10'h31c == io_inputs_0 ? 7'h0 : _GEN_3867; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3869 = 10'h31d == io_inputs_0 ? 7'h0 : _GEN_3868; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3870 = 10'h31e == io_inputs_0 ? 7'h0 : _GEN_3869; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3871 = 10'h31f == io_inputs_0 ? 7'h0 : _GEN_3870; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3872 = 10'h320 == io_inputs_0 ? 7'h0 : _GEN_3871; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3873 = 10'h321 == io_inputs_0 ? 7'h0 : _GEN_3872; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3874 = 10'h322 == io_inputs_0 ? 7'h0 : _GEN_3873; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3875 = 10'h323 == io_inputs_0 ? 7'h0 : _GEN_3874; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3876 = 10'h324 == io_inputs_0 ? 7'h0 : _GEN_3875; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3877 = 10'h325 == io_inputs_0 ? 7'h0 : _GEN_3876; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3878 = 10'h326 == io_inputs_0 ? 7'h0 : _GEN_3877; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3879 = 10'h327 == io_inputs_0 ? 7'h0 : _GEN_3878; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3880 = 10'h328 == io_inputs_0 ? 7'h0 : _GEN_3879; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3881 = 10'h329 == io_inputs_0 ? 7'h0 : _GEN_3880; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3882 = 10'h32a == io_inputs_0 ? 7'h0 : _GEN_3881; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3883 = 10'h32b == io_inputs_0 ? 7'h0 : _GEN_3882; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3884 = 10'h32c == io_inputs_0 ? 7'h0 : _GEN_3883; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3885 = 10'h32d == io_inputs_0 ? 7'h0 : _GEN_3884; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3886 = 10'h32e == io_inputs_0 ? 7'h0 : _GEN_3885; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3887 = 10'h32f == io_inputs_0 ? 7'h0 : _GEN_3886; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3888 = 10'h330 == io_inputs_0 ? 7'h0 : _GEN_3887; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3889 = 10'h331 == io_inputs_0 ? 7'h0 : _GEN_3888; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3890 = 10'h332 == io_inputs_0 ? 7'h0 : _GEN_3889; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3891 = 10'h333 == io_inputs_0 ? 7'h0 : _GEN_3890; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3892 = 10'h334 == io_inputs_0 ? 7'h0 : _GEN_3891; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3893 = 10'h335 == io_inputs_0 ? 7'h0 : _GEN_3892; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3894 = 10'h336 == io_inputs_0 ? 7'h0 : _GEN_3893; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3895 = 10'h337 == io_inputs_0 ? 7'h0 : _GEN_3894; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3896 = 10'h338 == io_inputs_0 ? 7'h0 : _GEN_3895; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3897 = 10'h339 == io_inputs_0 ? 7'h0 : _GEN_3896; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3898 = 10'h33a == io_inputs_0 ? 7'h0 : _GEN_3897; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3899 = 10'h33b == io_inputs_0 ? 7'h0 : _GEN_3898; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3900 = 10'h33c == io_inputs_0 ? 7'h0 : _GEN_3899; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3901 = 10'h33d == io_inputs_0 ? 7'h0 : _GEN_3900; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3902 = 10'h33e == io_inputs_0 ? 7'h0 : _GEN_3901; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3903 = 10'h33f == io_inputs_0 ? 7'h0 : _GEN_3902; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3904 = 10'h340 == io_inputs_0 ? 7'h0 : _GEN_3903; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3905 = 10'h341 == io_inputs_0 ? 7'h0 : _GEN_3904; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3906 = 10'h342 == io_inputs_0 ? 7'h0 : _GEN_3905; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3907 = 10'h343 == io_inputs_0 ? 7'h0 : _GEN_3906; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3908 = 10'h344 == io_inputs_0 ? 7'h0 : _GEN_3907; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3909 = 10'h345 == io_inputs_0 ? 7'h0 : _GEN_3908; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3910 = 10'h346 == io_inputs_0 ? 7'h0 : _GEN_3909; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3911 = 10'h347 == io_inputs_0 ? 7'h0 : _GEN_3910; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3912 = 10'h348 == io_inputs_0 ? 7'h0 : _GEN_3911; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3913 = 10'h349 == io_inputs_0 ? 7'h0 : _GEN_3912; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3914 = 10'h34a == io_inputs_0 ? 7'h0 : _GEN_3913; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3915 = 10'h34b == io_inputs_0 ? 7'h0 : _GEN_3914; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3916 = 10'h34c == io_inputs_0 ? 7'h0 : _GEN_3915; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3917 = 10'h34d == io_inputs_0 ? 7'h0 : _GEN_3916; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3918 = 10'h34e == io_inputs_0 ? 7'h0 : _GEN_3917; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3919 = 10'h34f == io_inputs_0 ? 7'h0 : _GEN_3918; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3920 = 10'h350 == io_inputs_0 ? 7'h0 : _GEN_3919; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3921 = 10'h351 == io_inputs_0 ? 7'h0 : _GEN_3920; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3922 = 10'h352 == io_inputs_0 ? 7'h0 : _GEN_3921; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3923 = 10'h353 == io_inputs_0 ? 7'h0 : _GEN_3922; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3924 = 10'h354 == io_inputs_0 ? 7'h0 : _GEN_3923; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3925 = 10'h355 == io_inputs_0 ? 7'h0 : _GEN_3924; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3926 = 10'h356 == io_inputs_0 ? 7'h0 : _GEN_3925; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3927 = 10'h357 == io_inputs_0 ? 7'h0 : _GEN_3926; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3928 = 10'h358 == io_inputs_0 ? 7'h0 : _GEN_3927; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3929 = 10'h359 == io_inputs_0 ? 7'h0 : _GEN_3928; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3930 = 10'h35a == io_inputs_0 ? 7'h0 : _GEN_3929; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3931 = 10'h35b == io_inputs_0 ? 7'h0 : _GEN_3930; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3932 = 10'h35c == io_inputs_0 ? 7'h0 : _GEN_3931; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3933 = 10'h35d == io_inputs_0 ? 7'h0 : _GEN_3932; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3934 = 10'h35e == io_inputs_0 ? 7'h0 : _GEN_3933; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3935 = 10'h35f == io_inputs_0 ? 7'h0 : _GEN_3934; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3936 = 10'h360 == io_inputs_0 ? 7'h0 : _GEN_3935; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3937 = 10'h361 == io_inputs_0 ? 7'h0 : _GEN_3936; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3938 = 10'h362 == io_inputs_0 ? 7'h0 : _GEN_3937; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3939 = 10'h363 == io_inputs_0 ? 7'h0 : _GEN_3938; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3940 = 10'h364 == io_inputs_0 ? 7'h0 : _GEN_3939; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3941 = 10'h365 == io_inputs_0 ? 7'h0 : _GEN_3940; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3942 = 10'h366 == io_inputs_0 ? 7'h0 : _GEN_3941; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3943 = 10'h367 == io_inputs_0 ? 7'h0 : _GEN_3942; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3944 = 10'h368 == io_inputs_0 ? 7'h0 : _GEN_3943; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3945 = 10'h369 == io_inputs_0 ? 7'h0 : _GEN_3944; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3946 = 10'h36a == io_inputs_0 ? 7'h0 : _GEN_3945; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3947 = 10'h36b == io_inputs_0 ? 7'h0 : _GEN_3946; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3948 = 10'h36c == io_inputs_0 ? 7'h0 : _GEN_3947; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3949 = 10'h36d == io_inputs_0 ? 7'h0 : _GEN_3948; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3950 = 10'h36e == io_inputs_0 ? 7'h0 : _GEN_3949; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3951 = 10'h36f == io_inputs_0 ? 7'h0 : _GEN_3950; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3952 = 10'h370 == io_inputs_0 ? 7'h0 : _GEN_3951; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3953 = 10'h371 == io_inputs_0 ? 7'h0 : _GEN_3952; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3954 = 10'h372 == io_inputs_0 ? 7'h0 : _GEN_3953; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3955 = 10'h373 == io_inputs_0 ? 7'h0 : _GEN_3954; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3956 = 10'h374 == io_inputs_0 ? 7'h0 : _GEN_3955; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3957 = 10'h375 == io_inputs_0 ? 7'h0 : _GEN_3956; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3958 = 10'h376 == io_inputs_0 ? 7'h0 : _GEN_3957; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3959 = 10'h377 == io_inputs_0 ? 7'h0 : _GEN_3958; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3960 = 10'h378 == io_inputs_0 ? 7'h0 : _GEN_3959; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3961 = 10'h379 == io_inputs_0 ? 7'h0 : _GEN_3960; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3962 = 10'h37a == io_inputs_0 ? 7'h0 : _GEN_3961; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3963 = 10'h37b == io_inputs_0 ? 7'h0 : _GEN_3962; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3964 = 10'h37c == io_inputs_0 ? 7'h0 : _GEN_3963; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3965 = 10'h37d == io_inputs_0 ? 7'h0 : _GEN_3964; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3966 = 10'h37e == io_inputs_0 ? 7'h0 : _GEN_3965; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3967 = 10'h37f == io_inputs_0 ? 7'h0 : _GEN_3966; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3968 = 10'h380 == io_inputs_0 ? 7'h0 : _GEN_3967; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3969 = 10'h381 == io_inputs_0 ? 7'h0 : _GEN_3968; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3970 = 10'h382 == io_inputs_0 ? 7'h0 : _GEN_3969; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3971 = 10'h383 == io_inputs_0 ? 7'h0 : _GEN_3970; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3972 = 10'h384 == io_inputs_0 ? 7'h0 : _GEN_3971; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3973 = 10'h385 == io_inputs_0 ? 7'h0 : _GEN_3972; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3974 = 10'h386 == io_inputs_0 ? 7'h0 : _GEN_3973; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3975 = 10'h387 == io_inputs_0 ? 7'h0 : _GEN_3974; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3976 = 10'h388 == io_inputs_0 ? 7'h0 : _GEN_3975; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3977 = 10'h389 == io_inputs_0 ? 7'h0 : _GEN_3976; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3978 = 10'h38a == io_inputs_0 ? 7'h0 : _GEN_3977; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3979 = 10'h38b == io_inputs_0 ? 7'h0 : _GEN_3978; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3980 = 10'h38c == io_inputs_0 ? 7'h0 : _GEN_3979; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3981 = 10'h38d == io_inputs_0 ? 7'h0 : _GEN_3980; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3982 = 10'h38e == io_inputs_0 ? 7'h0 : _GEN_3981; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3983 = 10'h38f == io_inputs_0 ? 7'h0 : _GEN_3982; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3984 = 10'h390 == io_inputs_0 ? 7'h0 : _GEN_3983; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3985 = 10'h391 == io_inputs_0 ? 7'h0 : _GEN_3984; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3986 = 10'h392 == io_inputs_0 ? 7'h0 : _GEN_3985; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3987 = 10'h393 == io_inputs_0 ? 7'h0 : _GEN_3986; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3988 = 10'h394 == io_inputs_0 ? 7'h0 : _GEN_3987; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3989 = 10'h395 == io_inputs_0 ? 7'h0 : _GEN_3988; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3990 = 10'h396 == io_inputs_0 ? 7'h0 : _GEN_3989; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3991 = 10'h397 == io_inputs_0 ? 7'h0 : _GEN_3990; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3992 = 10'h398 == io_inputs_0 ? 7'h0 : _GEN_3991; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3993 = 10'h399 == io_inputs_0 ? 7'h0 : _GEN_3992; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3994 = 10'h39a == io_inputs_0 ? 7'h0 : _GEN_3993; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3995 = 10'h39b == io_inputs_0 ? 7'h0 : _GEN_3994; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3996 = 10'h39c == io_inputs_0 ? 7'h0 : _GEN_3995; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3997 = 10'h39d == io_inputs_0 ? 7'h0 : _GEN_3996; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3998 = 10'h39e == io_inputs_0 ? 7'h0 : _GEN_3997; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_3999 = 10'h39f == io_inputs_0 ? 7'h0 : _GEN_3998; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4000 = 10'h3a0 == io_inputs_0 ? 7'h0 : _GEN_3999; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4001 = 10'h3a1 == io_inputs_0 ? 7'h0 : _GEN_4000; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4002 = 10'h3a2 == io_inputs_0 ? 7'h0 : _GEN_4001; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4003 = 10'h3a3 == io_inputs_0 ? 7'h0 : _GEN_4002; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4004 = 10'h3a4 == io_inputs_0 ? 7'h0 : _GEN_4003; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4005 = 10'h3a5 == io_inputs_0 ? 7'h0 : _GEN_4004; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4006 = 10'h3a6 == io_inputs_0 ? 7'h0 : _GEN_4005; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4007 = 10'h3a7 == io_inputs_0 ? 7'h0 : _GEN_4006; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4008 = 10'h3a8 == io_inputs_0 ? 7'h0 : _GEN_4007; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4009 = 10'h3a9 == io_inputs_0 ? 7'h0 : _GEN_4008; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4010 = 10'h3aa == io_inputs_0 ? 7'h0 : _GEN_4009; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4011 = 10'h3ab == io_inputs_0 ? 7'h0 : _GEN_4010; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4012 = 10'h3ac == io_inputs_0 ? 7'h0 : _GEN_4011; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4013 = 10'h3ad == io_inputs_0 ? 7'h0 : _GEN_4012; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4014 = 10'h3ae == io_inputs_0 ? 7'h0 : _GEN_4013; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4015 = 10'h3af == io_inputs_0 ? 7'h0 : _GEN_4014; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4016 = 10'h3b0 == io_inputs_0 ? 7'h0 : _GEN_4015; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4017 = 10'h3b1 == io_inputs_0 ? 7'h0 : _GEN_4016; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4018 = 10'h3b2 == io_inputs_0 ? 7'h0 : _GEN_4017; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4019 = 10'h3b3 == io_inputs_0 ? 7'h0 : _GEN_4018; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4020 = 10'h3b4 == io_inputs_0 ? 7'h0 : _GEN_4019; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4021 = 10'h3b5 == io_inputs_0 ? 7'h0 : _GEN_4020; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4022 = 10'h3b6 == io_inputs_0 ? 7'h0 : _GEN_4021; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4023 = 10'h3b7 == io_inputs_0 ? 7'h0 : _GEN_4022; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4024 = 10'h3b8 == io_inputs_0 ? 7'h0 : _GEN_4023; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4025 = 10'h3b9 == io_inputs_0 ? 7'h0 : _GEN_4024; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4026 = 10'h3ba == io_inputs_0 ? 7'h0 : _GEN_4025; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4027 = 10'h3bb == io_inputs_0 ? 7'h0 : _GEN_4026; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4028 = 10'h3bc == io_inputs_0 ? 7'h0 : _GEN_4027; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4029 = 10'h3bd == io_inputs_0 ? 7'h0 : _GEN_4028; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4030 = 10'h3be == io_inputs_0 ? 7'h0 : _GEN_4029; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4031 = 10'h3bf == io_inputs_0 ? 7'h0 : _GEN_4030; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4032 = 10'h3c0 == io_inputs_0 ? 7'h0 : _GEN_4031; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4033 = 10'h3c1 == io_inputs_0 ? 7'h0 : _GEN_4032; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4034 = 10'h3c2 == io_inputs_0 ? 7'h0 : _GEN_4033; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4035 = 10'h3c3 == io_inputs_0 ? 7'h0 : _GEN_4034; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4036 = 10'h3c4 == io_inputs_0 ? 7'h0 : _GEN_4035; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4037 = 10'h3c5 == io_inputs_0 ? 7'h0 : _GEN_4036; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4038 = 10'h3c6 == io_inputs_0 ? 7'h0 : _GEN_4037; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4039 = 10'h3c7 == io_inputs_0 ? 7'h0 : _GEN_4038; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4040 = 10'h3c8 == io_inputs_0 ? 7'h0 : _GEN_4039; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4041 = 10'h3c9 == io_inputs_0 ? 7'h0 : _GEN_4040; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4042 = 10'h3ca == io_inputs_0 ? 7'h0 : _GEN_4041; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4043 = 10'h3cb == io_inputs_0 ? 7'h0 : _GEN_4042; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4044 = 10'h3cc == io_inputs_0 ? 7'h0 : _GEN_4043; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4045 = 10'h3cd == io_inputs_0 ? 7'h0 : _GEN_4044; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4046 = 10'h3ce == io_inputs_0 ? 7'h0 : _GEN_4045; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4047 = 10'h3cf == io_inputs_0 ? 7'h0 : _GEN_4046; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4048 = 10'h3d0 == io_inputs_0 ? 7'h0 : _GEN_4047; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4049 = 10'h3d1 == io_inputs_0 ? 7'h0 : _GEN_4048; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4050 = 10'h3d2 == io_inputs_0 ? 7'h0 : _GEN_4049; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4051 = 10'h3d3 == io_inputs_0 ? 7'h0 : _GEN_4050; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4052 = 10'h3d4 == io_inputs_0 ? 7'h0 : _GEN_4051; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4053 = 10'h3d5 == io_inputs_0 ? 7'h0 : _GEN_4052; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4054 = 10'h3d6 == io_inputs_0 ? 7'h0 : _GEN_4053; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4055 = 10'h3d7 == io_inputs_0 ? 7'h0 : _GEN_4054; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4056 = 10'h3d8 == io_inputs_0 ? 7'h0 : _GEN_4055; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4057 = 10'h3d9 == io_inputs_0 ? 7'h0 : _GEN_4056; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4058 = 10'h3da == io_inputs_0 ? 7'h0 : _GEN_4057; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4059 = 10'h3db == io_inputs_0 ? 7'h0 : _GEN_4058; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4060 = 10'h3dc == io_inputs_0 ? 7'h0 : _GEN_4059; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4061 = 10'h3dd == io_inputs_0 ? 7'h0 : _GEN_4060; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4062 = 10'h3de == io_inputs_0 ? 7'h0 : _GEN_4061; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4063 = 10'h3df == io_inputs_0 ? 7'h0 : _GEN_4062; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4064 = 10'h3e0 == io_inputs_0 ? 7'h0 : _GEN_4063; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4065 = 10'h3e1 == io_inputs_0 ? 7'h0 : _GEN_4064; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4066 = 10'h3e2 == io_inputs_0 ? 7'h0 : _GEN_4065; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4067 = 10'h3e3 == io_inputs_0 ? 7'h0 : _GEN_4066; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4068 = 10'h3e4 == io_inputs_0 ? 7'h0 : _GEN_4067; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4069 = 10'h3e5 == io_inputs_0 ? 7'h0 : _GEN_4068; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4070 = 10'h3e6 == io_inputs_0 ? 7'h0 : _GEN_4069; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4071 = 10'h3e7 == io_inputs_0 ? 7'h0 : _GEN_4070; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4072 = 10'h3e8 == io_inputs_0 ? 7'h0 : _GEN_4071; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4073 = 10'h3e9 == io_inputs_0 ? 7'h0 : _GEN_4072; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4074 = 10'h3ea == io_inputs_0 ? 7'h0 : _GEN_4073; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4075 = 10'h3eb == io_inputs_0 ? 7'h0 : _GEN_4074; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4076 = 10'h3ec == io_inputs_0 ? 7'h0 : _GEN_4075; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4077 = 10'h3ed == io_inputs_0 ? 7'h0 : _GEN_4076; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4078 = 10'h3ee == io_inputs_0 ? 7'h0 : _GEN_4077; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4079 = 10'h3ef == io_inputs_0 ? 7'h0 : _GEN_4078; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4080 = 10'h3f0 == io_inputs_0 ? 7'h0 : _GEN_4079; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4081 = 10'h3f1 == io_inputs_0 ? 7'h0 : _GEN_4080; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4082 = 10'h3f2 == io_inputs_0 ? 7'h0 : _GEN_4081; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4083 = 10'h3f3 == io_inputs_0 ? 7'h0 : _GEN_4082; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4084 = 10'h3f4 == io_inputs_0 ? 7'h0 : _GEN_4083; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4085 = 10'h3f5 == io_inputs_0 ? 7'h0 : _GEN_4084; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4086 = 10'h3f6 == io_inputs_0 ? 7'h0 : _GEN_4085; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4087 = 10'h3f7 == io_inputs_0 ? 7'h0 : _GEN_4086; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4088 = 10'h3f8 == io_inputs_0 ? 7'h0 : _GEN_4087; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4089 = 10'h3f9 == io_inputs_0 ? 7'h0 : _GEN_4088; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4090 = 10'h3fa == io_inputs_0 ? 7'h0 : _GEN_4089; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4091 = 10'h3fb == io_inputs_0 ? 7'h0 : _GEN_4090; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4092 = 10'h3fc == io_inputs_0 ? 7'h0 : _GEN_4091; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4597 = 10'h1f5 == io_inputs_0 ? 7'h1 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4598 = 10'h1f6 == io_inputs_0 ? 7'h2 : _GEN_4597; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4599 = 10'h1f7 == io_inputs_0 ? 7'h3 : _GEN_4598; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4600 = 10'h1f8 == io_inputs_0 ? 7'h4 : _GEN_4599; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4601 = 10'h1f9 == io_inputs_0 ? 7'h5 : _GEN_4600; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4602 = 10'h1fa == io_inputs_0 ? 7'h6 : _GEN_4601; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4603 = 10'h1fb == io_inputs_0 ? 7'h7 : _GEN_4602; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4604 = 10'h1fc == io_inputs_0 ? 7'h8 : _GEN_4603; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4605 = 10'h1fd == io_inputs_0 ? 7'h9 : _GEN_4604; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4606 = 10'h1fe == io_inputs_0 ? 7'ha : _GEN_4605; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4607 = 10'h1ff == io_inputs_0 ? 7'hb : _GEN_4606; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4608 = 10'h200 == io_inputs_0 ? 7'hc : _GEN_4607; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4609 = 10'h201 == io_inputs_0 ? 7'hd : _GEN_4608; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4610 = 10'h202 == io_inputs_0 ? 7'he : _GEN_4609; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4611 = 10'h203 == io_inputs_0 ? 7'hf : _GEN_4610; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4612 = 10'h204 == io_inputs_0 ? 7'h10 : _GEN_4611; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4613 = 10'h205 == io_inputs_0 ? 7'h11 : _GEN_4612; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4614 = 10'h206 == io_inputs_0 ? 7'h12 : _GEN_4613; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4615 = 10'h207 == io_inputs_0 ? 7'h13 : _GEN_4614; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4616 = 10'h208 == io_inputs_0 ? 7'h14 : _GEN_4615; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4617 = 10'h209 == io_inputs_0 ? 7'h15 : _GEN_4616; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4618 = 10'h20a == io_inputs_0 ? 7'h16 : _GEN_4617; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4619 = 10'h20b == io_inputs_0 ? 7'h17 : _GEN_4618; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4620 = 10'h20c == io_inputs_0 ? 7'h18 : _GEN_4619; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4621 = 10'h20d == io_inputs_0 ? 7'h19 : _GEN_4620; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4622 = 10'h20e == io_inputs_0 ? 7'h1a : _GEN_4621; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4623 = 10'h20f == io_inputs_0 ? 7'h1b : _GEN_4622; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4624 = 10'h210 == io_inputs_0 ? 7'h1c : _GEN_4623; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4625 = 10'h211 == io_inputs_0 ? 7'h1d : _GEN_4624; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4626 = 10'h212 == io_inputs_0 ? 7'h1e : _GEN_4625; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4627 = 10'h213 == io_inputs_0 ? 7'h1f : _GEN_4626; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4628 = 10'h214 == io_inputs_0 ? 7'h20 : _GEN_4627; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4629 = 10'h215 == io_inputs_0 ? 7'h21 : _GEN_4628; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4630 = 10'h216 == io_inputs_0 ? 7'h22 : _GEN_4629; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4631 = 10'h217 == io_inputs_0 ? 7'h23 : _GEN_4630; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4632 = 10'h218 == io_inputs_0 ? 7'h24 : _GEN_4631; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4633 = 10'h219 == io_inputs_0 ? 7'h25 : _GEN_4632; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4634 = 10'h21a == io_inputs_0 ? 7'h26 : _GEN_4633; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4635 = 10'h21b == io_inputs_0 ? 7'h27 : _GEN_4634; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4636 = 10'h21c == io_inputs_0 ? 7'h28 : _GEN_4635; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4637 = 10'h21d == io_inputs_0 ? 7'h29 : _GEN_4636; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4638 = 10'h21e == io_inputs_0 ? 7'h2a : _GEN_4637; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4639 = 10'h21f == io_inputs_0 ? 7'h2b : _GEN_4638; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4640 = 10'h220 == io_inputs_0 ? 7'h2c : _GEN_4639; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4641 = 10'h221 == io_inputs_0 ? 7'h2d : _GEN_4640; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4642 = 10'h222 == io_inputs_0 ? 7'h2e : _GEN_4641; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4643 = 10'h223 == io_inputs_0 ? 7'h2f : _GEN_4642; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4644 = 10'h224 == io_inputs_0 ? 7'h30 : _GEN_4643; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4645 = 10'h225 == io_inputs_0 ? 7'h31 : _GEN_4644; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4646 = 10'h226 == io_inputs_0 ? 7'h32 : _GEN_4645; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4647 = 10'h227 == io_inputs_0 ? 7'h33 : _GEN_4646; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4648 = 10'h228 == io_inputs_0 ? 7'h34 : _GEN_4647; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4649 = 10'h229 == io_inputs_0 ? 7'h35 : _GEN_4648; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4650 = 10'h22a == io_inputs_0 ? 7'h36 : _GEN_4649; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4651 = 10'h22b == io_inputs_0 ? 7'h37 : _GEN_4650; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4652 = 10'h22c == io_inputs_0 ? 7'h38 : _GEN_4651; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4653 = 10'h22d == io_inputs_0 ? 7'h39 : _GEN_4652; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4654 = 10'h22e == io_inputs_0 ? 7'h3a : _GEN_4653; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4655 = 10'h22f == io_inputs_0 ? 7'h3b : _GEN_4654; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4656 = 10'h230 == io_inputs_0 ? 7'h3c : _GEN_4655; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4657 = 10'h231 == io_inputs_0 ? 7'h3d : _GEN_4656; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4658 = 10'h232 == io_inputs_0 ? 7'h3e : _GEN_4657; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4659 = 10'h233 == io_inputs_0 ? 7'h3f : _GEN_4658; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4660 = 10'h234 == io_inputs_0 ? 7'h40 : _GEN_4659; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4661 = 10'h235 == io_inputs_0 ? 7'h41 : _GEN_4660; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4662 = 10'h236 == io_inputs_0 ? 7'h42 : _GEN_4661; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4663 = 10'h237 == io_inputs_0 ? 7'h43 : _GEN_4662; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4664 = 10'h238 == io_inputs_0 ? 7'h44 : _GEN_4663; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4665 = 10'h239 == io_inputs_0 ? 7'h45 : _GEN_4664; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4666 = 10'h23a == io_inputs_0 ? 7'h46 : _GEN_4665; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4667 = 10'h23b == io_inputs_0 ? 7'h47 : _GEN_4666; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4668 = 10'h23c == io_inputs_0 ? 7'h48 : _GEN_4667; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4669 = 10'h23d == io_inputs_0 ? 7'h49 : _GEN_4668; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4670 = 10'h23e == io_inputs_0 ? 7'h4a : _GEN_4669; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4671 = 10'h23f == io_inputs_0 ? 7'h4b : _GEN_4670; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4672 = 10'h240 == io_inputs_0 ? 7'h4c : _GEN_4671; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4673 = 10'h241 == io_inputs_0 ? 7'h4d : _GEN_4672; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4674 = 10'h242 == io_inputs_0 ? 7'h4e : _GEN_4673; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4675 = 10'h243 == io_inputs_0 ? 7'h4f : _GEN_4674; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4676 = 10'h244 == io_inputs_0 ? 7'h50 : _GEN_4675; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4677 = 10'h245 == io_inputs_0 ? 7'h51 : _GEN_4676; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4678 = 10'h246 == io_inputs_0 ? 7'h52 : _GEN_4677; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4679 = 10'h247 == io_inputs_0 ? 7'h53 : _GEN_4678; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4680 = 10'h248 == io_inputs_0 ? 7'h54 : _GEN_4679; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4681 = 10'h249 == io_inputs_0 ? 7'h55 : _GEN_4680; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4682 = 10'h24a == io_inputs_0 ? 7'h56 : _GEN_4681; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4683 = 10'h24b == io_inputs_0 ? 7'h57 : _GEN_4682; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4684 = 10'h24c == io_inputs_0 ? 7'h58 : _GEN_4683; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4685 = 10'h24d == io_inputs_0 ? 7'h59 : _GEN_4684; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4686 = 10'h24e == io_inputs_0 ? 7'h5a : _GEN_4685; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4687 = 10'h24f == io_inputs_0 ? 7'h5b : _GEN_4686; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4688 = 10'h250 == io_inputs_0 ? 7'h5c : _GEN_4687; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4689 = 10'h251 == io_inputs_0 ? 7'h5d : _GEN_4688; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4690 = 10'h252 == io_inputs_0 ? 7'h5e : _GEN_4689; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4691 = 10'h253 == io_inputs_0 ? 7'h5f : _GEN_4690; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4692 = 10'h254 == io_inputs_0 ? 7'h60 : _GEN_4691; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4693 = 10'h255 == io_inputs_0 ? 7'h61 : _GEN_4692; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4694 = 10'h256 == io_inputs_0 ? 7'h62 : _GEN_4693; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4695 = 10'h257 == io_inputs_0 ? 7'h63 : _GEN_4694; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4696 = 10'h258 == io_inputs_0 ? 7'h64 : _GEN_4695; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4697 = 10'h259 == io_inputs_0 ? 7'h64 : _GEN_4696; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4698 = 10'h25a == io_inputs_0 ? 7'h64 : _GEN_4697; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4699 = 10'h25b == io_inputs_0 ? 7'h64 : _GEN_4698; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4700 = 10'h25c == io_inputs_0 ? 7'h64 : _GEN_4699; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4701 = 10'h25d == io_inputs_0 ? 7'h64 : _GEN_4700; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4702 = 10'h25e == io_inputs_0 ? 7'h64 : _GEN_4701; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4703 = 10'h25f == io_inputs_0 ? 7'h64 : _GEN_4702; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4704 = 10'h260 == io_inputs_0 ? 7'h64 : _GEN_4703; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4705 = 10'h261 == io_inputs_0 ? 7'h64 : _GEN_4704; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4706 = 10'h262 == io_inputs_0 ? 7'h64 : _GEN_4705; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4707 = 10'h263 == io_inputs_0 ? 7'h64 : _GEN_4706; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4708 = 10'h264 == io_inputs_0 ? 7'h64 : _GEN_4707; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4709 = 10'h265 == io_inputs_0 ? 7'h64 : _GEN_4708; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4710 = 10'h266 == io_inputs_0 ? 7'h64 : _GEN_4709; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4711 = 10'h267 == io_inputs_0 ? 7'h64 : _GEN_4710; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4712 = 10'h268 == io_inputs_0 ? 7'h64 : _GEN_4711; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4713 = 10'h269 == io_inputs_0 ? 7'h64 : _GEN_4712; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4714 = 10'h26a == io_inputs_0 ? 7'h64 : _GEN_4713; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4715 = 10'h26b == io_inputs_0 ? 7'h64 : _GEN_4714; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4716 = 10'h26c == io_inputs_0 ? 7'h64 : _GEN_4715; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4717 = 10'h26d == io_inputs_0 ? 7'h64 : _GEN_4716; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4718 = 10'h26e == io_inputs_0 ? 7'h64 : _GEN_4717; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4719 = 10'h26f == io_inputs_0 ? 7'h64 : _GEN_4718; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4720 = 10'h270 == io_inputs_0 ? 7'h64 : _GEN_4719; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4721 = 10'h271 == io_inputs_0 ? 7'h64 : _GEN_4720; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4722 = 10'h272 == io_inputs_0 ? 7'h64 : _GEN_4721; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4723 = 10'h273 == io_inputs_0 ? 7'h64 : _GEN_4722; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4724 = 10'h274 == io_inputs_0 ? 7'h64 : _GEN_4723; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4725 = 10'h275 == io_inputs_0 ? 7'h64 : _GEN_4724; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4726 = 10'h276 == io_inputs_0 ? 7'h64 : _GEN_4725; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4727 = 10'h277 == io_inputs_0 ? 7'h64 : _GEN_4726; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4728 = 10'h278 == io_inputs_0 ? 7'h64 : _GEN_4727; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4729 = 10'h279 == io_inputs_0 ? 7'h64 : _GEN_4728; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4730 = 10'h27a == io_inputs_0 ? 7'h64 : _GEN_4729; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4731 = 10'h27b == io_inputs_0 ? 7'h64 : _GEN_4730; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4732 = 10'h27c == io_inputs_0 ? 7'h64 : _GEN_4731; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4733 = 10'h27d == io_inputs_0 ? 7'h64 : _GEN_4732; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4734 = 10'h27e == io_inputs_0 ? 7'h64 : _GEN_4733; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4735 = 10'h27f == io_inputs_0 ? 7'h64 : _GEN_4734; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4736 = 10'h280 == io_inputs_0 ? 7'h64 : _GEN_4735; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4737 = 10'h281 == io_inputs_0 ? 7'h64 : _GEN_4736; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4738 = 10'h282 == io_inputs_0 ? 7'h64 : _GEN_4737; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4739 = 10'h283 == io_inputs_0 ? 7'h64 : _GEN_4738; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4740 = 10'h284 == io_inputs_0 ? 7'h64 : _GEN_4739; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4741 = 10'h285 == io_inputs_0 ? 7'h64 : _GEN_4740; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4742 = 10'h286 == io_inputs_0 ? 7'h64 : _GEN_4741; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4743 = 10'h287 == io_inputs_0 ? 7'h64 : _GEN_4742; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4744 = 10'h288 == io_inputs_0 ? 7'h64 : _GEN_4743; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4745 = 10'h289 == io_inputs_0 ? 7'h64 : _GEN_4744; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4746 = 10'h28a == io_inputs_0 ? 7'h64 : _GEN_4745; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4747 = 10'h28b == io_inputs_0 ? 7'h64 : _GEN_4746; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4748 = 10'h28c == io_inputs_0 ? 7'h64 : _GEN_4747; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4749 = 10'h28d == io_inputs_0 ? 7'h64 : _GEN_4748; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4750 = 10'h28e == io_inputs_0 ? 7'h64 : _GEN_4749; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4751 = 10'h28f == io_inputs_0 ? 7'h64 : _GEN_4750; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4752 = 10'h290 == io_inputs_0 ? 7'h64 : _GEN_4751; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4753 = 10'h291 == io_inputs_0 ? 7'h64 : _GEN_4752; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4754 = 10'h292 == io_inputs_0 ? 7'h64 : _GEN_4753; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4755 = 10'h293 == io_inputs_0 ? 7'h64 : _GEN_4754; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4756 = 10'h294 == io_inputs_0 ? 7'h64 : _GEN_4755; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4757 = 10'h295 == io_inputs_0 ? 7'h64 : _GEN_4756; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4758 = 10'h296 == io_inputs_0 ? 7'h64 : _GEN_4757; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4759 = 10'h297 == io_inputs_0 ? 7'h64 : _GEN_4758; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4760 = 10'h298 == io_inputs_0 ? 7'h64 : _GEN_4759; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4761 = 10'h299 == io_inputs_0 ? 7'h64 : _GEN_4760; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4762 = 10'h29a == io_inputs_0 ? 7'h64 : _GEN_4761; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4763 = 10'h29b == io_inputs_0 ? 7'h64 : _GEN_4762; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4764 = 10'h29c == io_inputs_0 ? 7'h64 : _GEN_4763; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4765 = 10'h29d == io_inputs_0 ? 7'h64 : _GEN_4764; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4766 = 10'h29e == io_inputs_0 ? 7'h64 : _GEN_4765; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4767 = 10'h29f == io_inputs_0 ? 7'h64 : _GEN_4766; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4768 = 10'h2a0 == io_inputs_0 ? 7'h64 : _GEN_4767; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4769 = 10'h2a1 == io_inputs_0 ? 7'h64 : _GEN_4768; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4770 = 10'h2a2 == io_inputs_0 ? 7'h64 : _GEN_4769; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4771 = 10'h2a3 == io_inputs_0 ? 7'h64 : _GEN_4770; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4772 = 10'h2a4 == io_inputs_0 ? 7'h64 : _GEN_4771; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4773 = 10'h2a5 == io_inputs_0 ? 7'h64 : _GEN_4772; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4774 = 10'h2a6 == io_inputs_0 ? 7'h64 : _GEN_4773; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4775 = 10'h2a7 == io_inputs_0 ? 7'h64 : _GEN_4774; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4776 = 10'h2a8 == io_inputs_0 ? 7'h64 : _GEN_4775; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4777 = 10'h2a9 == io_inputs_0 ? 7'h64 : _GEN_4776; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4778 = 10'h2aa == io_inputs_0 ? 7'h64 : _GEN_4777; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4779 = 10'h2ab == io_inputs_0 ? 7'h64 : _GEN_4778; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4780 = 10'h2ac == io_inputs_0 ? 7'h64 : _GEN_4779; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4781 = 10'h2ad == io_inputs_0 ? 7'h64 : _GEN_4780; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4782 = 10'h2ae == io_inputs_0 ? 7'h64 : _GEN_4781; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4783 = 10'h2af == io_inputs_0 ? 7'h64 : _GEN_4782; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4784 = 10'h2b0 == io_inputs_0 ? 7'h64 : _GEN_4783; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4785 = 10'h2b1 == io_inputs_0 ? 7'h64 : _GEN_4784; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4786 = 10'h2b2 == io_inputs_0 ? 7'h64 : _GEN_4785; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4787 = 10'h2b3 == io_inputs_0 ? 7'h64 : _GEN_4786; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4788 = 10'h2b4 == io_inputs_0 ? 7'h64 : _GEN_4787; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4789 = 10'h2b5 == io_inputs_0 ? 7'h64 : _GEN_4788; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4790 = 10'h2b6 == io_inputs_0 ? 7'h64 : _GEN_4789; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4791 = 10'h2b7 == io_inputs_0 ? 7'h64 : _GEN_4790; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4792 = 10'h2b8 == io_inputs_0 ? 7'h64 : _GEN_4791; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4793 = 10'h2b9 == io_inputs_0 ? 7'h64 : _GEN_4792; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4794 = 10'h2ba == io_inputs_0 ? 7'h64 : _GEN_4793; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4795 = 10'h2bb == io_inputs_0 ? 7'h64 : _GEN_4794; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4796 = 10'h2bc == io_inputs_0 ? 7'h64 : _GEN_4795; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4797 = 10'h2bd == io_inputs_0 ? 7'h64 : _GEN_4796; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4798 = 10'h2be == io_inputs_0 ? 7'h64 : _GEN_4797; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4799 = 10'h2bf == io_inputs_0 ? 7'h64 : _GEN_4798; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4800 = 10'h2c0 == io_inputs_0 ? 7'h64 : _GEN_4799; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4801 = 10'h2c1 == io_inputs_0 ? 7'h64 : _GEN_4800; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4802 = 10'h2c2 == io_inputs_0 ? 7'h64 : _GEN_4801; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4803 = 10'h2c3 == io_inputs_0 ? 7'h64 : _GEN_4802; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4804 = 10'h2c4 == io_inputs_0 ? 7'h64 : _GEN_4803; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4805 = 10'h2c5 == io_inputs_0 ? 7'h64 : _GEN_4804; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4806 = 10'h2c6 == io_inputs_0 ? 7'h64 : _GEN_4805; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4807 = 10'h2c7 == io_inputs_0 ? 7'h64 : _GEN_4806; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4808 = 10'h2c8 == io_inputs_0 ? 7'h64 : _GEN_4807; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4809 = 10'h2c9 == io_inputs_0 ? 7'h64 : _GEN_4808; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4810 = 10'h2ca == io_inputs_0 ? 7'h64 : _GEN_4809; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4811 = 10'h2cb == io_inputs_0 ? 7'h64 : _GEN_4810; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4812 = 10'h2cc == io_inputs_0 ? 7'h64 : _GEN_4811; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4813 = 10'h2cd == io_inputs_0 ? 7'h64 : _GEN_4812; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4814 = 10'h2ce == io_inputs_0 ? 7'h64 : _GEN_4813; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4815 = 10'h2cf == io_inputs_0 ? 7'h64 : _GEN_4814; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4816 = 10'h2d0 == io_inputs_0 ? 7'h64 : _GEN_4815; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4817 = 10'h2d1 == io_inputs_0 ? 7'h64 : _GEN_4816; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4818 = 10'h2d2 == io_inputs_0 ? 7'h64 : _GEN_4817; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4819 = 10'h2d3 == io_inputs_0 ? 7'h64 : _GEN_4818; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4820 = 10'h2d4 == io_inputs_0 ? 7'h64 : _GEN_4819; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4821 = 10'h2d5 == io_inputs_0 ? 7'h64 : _GEN_4820; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4822 = 10'h2d6 == io_inputs_0 ? 7'h64 : _GEN_4821; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4823 = 10'h2d7 == io_inputs_0 ? 7'h64 : _GEN_4822; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4824 = 10'h2d8 == io_inputs_0 ? 7'h64 : _GEN_4823; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4825 = 10'h2d9 == io_inputs_0 ? 7'h64 : _GEN_4824; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4826 = 10'h2da == io_inputs_0 ? 7'h64 : _GEN_4825; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4827 = 10'h2db == io_inputs_0 ? 7'h64 : _GEN_4826; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4828 = 10'h2dc == io_inputs_0 ? 7'h64 : _GEN_4827; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4829 = 10'h2dd == io_inputs_0 ? 7'h64 : _GEN_4828; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4830 = 10'h2de == io_inputs_0 ? 7'h64 : _GEN_4829; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4831 = 10'h2df == io_inputs_0 ? 7'h64 : _GEN_4830; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4832 = 10'h2e0 == io_inputs_0 ? 7'h64 : _GEN_4831; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4833 = 10'h2e1 == io_inputs_0 ? 7'h64 : _GEN_4832; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4834 = 10'h2e2 == io_inputs_0 ? 7'h64 : _GEN_4833; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4835 = 10'h2e3 == io_inputs_0 ? 7'h64 : _GEN_4834; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4836 = 10'h2e4 == io_inputs_0 ? 7'h64 : _GEN_4835; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4837 = 10'h2e5 == io_inputs_0 ? 7'h64 : _GEN_4836; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4838 = 10'h2e6 == io_inputs_0 ? 7'h64 : _GEN_4837; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4839 = 10'h2e7 == io_inputs_0 ? 7'h64 : _GEN_4838; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4840 = 10'h2e8 == io_inputs_0 ? 7'h64 : _GEN_4839; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4841 = 10'h2e9 == io_inputs_0 ? 7'h64 : _GEN_4840; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4842 = 10'h2ea == io_inputs_0 ? 7'h64 : _GEN_4841; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4843 = 10'h2eb == io_inputs_0 ? 7'h64 : _GEN_4842; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4844 = 10'h2ec == io_inputs_0 ? 7'h64 : _GEN_4843; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4845 = 10'h2ed == io_inputs_0 ? 7'h64 : _GEN_4844; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4846 = 10'h2ee == io_inputs_0 ? 7'h64 : _GEN_4845; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4847 = 10'h2ef == io_inputs_0 ? 7'h64 : _GEN_4846; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4848 = 10'h2f0 == io_inputs_0 ? 7'h64 : _GEN_4847; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4849 = 10'h2f1 == io_inputs_0 ? 7'h64 : _GEN_4848; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4850 = 10'h2f2 == io_inputs_0 ? 7'h64 : _GEN_4849; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4851 = 10'h2f3 == io_inputs_0 ? 7'h64 : _GEN_4850; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4852 = 10'h2f4 == io_inputs_0 ? 7'h64 : _GEN_4851; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4853 = 10'h2f5 == io_inputs_0 ? 7'h64 : _GEN_4852; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4854 = 10'h2f6 == io_inputs_0 ? 7'h64 : _GEN_4853; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4855 = 10'h2f7 == io_inputs_0 ? 7'h64 : _GEN_4854; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4856 = 10'h2f8 == io_inputs_0 ? 7'h64 : _GEN_4855; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4857 = 10'h2f9 == io_inputs_0 ? 7'h64 : _GEN_4856; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4858 = 10'h2fa == io_inputs_0 ? 7'h64 : _GEN_4857; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4859 = 10'h2fb == io_inputs_0 ? 7'h64 : _GEN_4858; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4860 = 10'h2fc == io_inputs_0 ? 7'h64 : _GEN_4859; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4861 = 10'h2fd == io_inputs_0 ? 7'h64 : _GEN_4860; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4862 = 10'h2fe == io_inputs_0 ? 7'h64 : _GEN_4861; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4863 = 10'h2ff == io_inputs_0 ? 7'h64 : _GEN_4862; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4864 = 10'h300 == io_inputs_0 ? 7'h64 : _GEN_4863; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4865 = 10'h301 == io_inputs_0 ? 7'h64 : _GEN_4864; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4866 = 10'h302 == io_inputs_0 ? 7'h64 : _GEN_4865; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4867 = 10'h303 == io_inputs_0 ? 7'h64 : _GEN_4866; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4868 = 10'h304 == io_inputs_0 ? 7'h64 : _GEN_4867; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4869 = 10'h305 == io_inputs_0 ? 7'h64 : _GEN_4868; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4870 = 10'h306 == io_inputs_0 ? 7'h64 : _GEN_4869; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4871 = 10'h307 == io_inputs_0 ? 7'h64 : _GEN_4870; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4872 = 10'h308 == io_inputs_0 ? 7'h64 : _GEN_4871; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4873 = 10'h309 == io_inputs_0 ? 7'h64 : _GEN_4872; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4874 = 10'h30a == io_inputs_0 ? 7'h64 : _GEN_4873; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4875 = 10'h30b == io_inputs_0 ? 7'h64 : _GEN_4874; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4876 = 10'h30c == io_inputs_0 ? 7'h64 : _GEN_4875; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4877 = 10'h30d == io_inputs_0 ? 7'h64 : _GEN_4876; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4878 = 10'h30e == io_inputs_0 ? 7'h64 : _GEN_4877; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4879 = 10'h30f == io_inputs_0 ? 7'h64 : _GEN_4878; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4880 = 10'h310 == io_inputs_0 ? 7'h64 : _GEN_4879; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4881 = 10'h311 == io_inputs_0 ? 7'h64 : _GEN_4880; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4882 = 10'h312 == io_inputs_0 ? 7'h64 : _GEN_4881; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4883 = 10'h313 == io_inputs_0 ? 7'h64 : _GEN_4882; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4884 = 10'h314 == io_inputs_0 ? 7'h64 : _GEN_4883; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4885 = 10'h315 == io_inputs_0 ? 7'h64 : _GEN_4884; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4886 = 10'h316 == io_inputs_0 ? 7'h64 : _GEN_4885; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4887 = 10'h317 == io_inputs_0 ? 7'h64 : _GEN_4886; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4888 = 10'h318 == io_inputs_0 ? 7'h64 : _GEN_4887; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4889 = 10'h319 == io_inputs_0 ? 7'h64 : _GEN_4888; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4890 = 10'h31a == io_inputs_0 ? 7'h64 : _GEN_4889; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4891 = 10'h31b == io_inputs_0 ? 7'h64 : _GEN_4890; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4892 = 10'h31c == io_inputs_0 ? 7'h64 : _GEN_4891; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4893 = 10'h31d == io_inputs_0 ? 7'h64 : _GEN_4892; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4894 = 10'h31e == io_inputs_0 ? 7'h64 : _GEN_4893; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4895 = 10'h31f == io_inputs_0 ? 7'h64 : _GEN_4894; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4896 = 10'h320 == io_inputs_0 ? 7'h64 : _GEN_4895; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4897 = 10'h321 == io_inputs_0 ? 7'h64 : _GEN_4896; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4898 = 10'h322 == io_inputs_0 ? 7'h64 : _GEN_4897; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4899 = 10'h323 == io_inputs_0 ? 7'h64 : _GEN_4898; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4900 = 10'h324 == io_inputs_0 ? 7'h64 : _GEN_4899; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4901 = 10'h325 == io_inputs_0 ? 7'h64 : _GEN_4900; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4902 = 10'h326 == io_inputs_0 ? 7'h64 : _GEN_4901; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4903 = 10'h327 == io_inputs_0 ? 7'h64 : _GEN_4902; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4904 = 10'h328 == io_inputs_0 ? 7'h64 : _GEN_4903; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4905 = 10'h329 == io_inputs_0 ? 7'h64 : _GEN_4904; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4906 = 10'h32a == io_inputs_0 ? 7'h64 : _GEN_4905; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4907 = 10'h32b == io_inputs_0 ? 7'h64 : _GEN_4906; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4908 = 10'h32c == io_inputs_0 ? 7'h64 : _GEN_4907; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4909 = 10'h32d == io_inputs_0 ? 7'h64 : _GEN_4908; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4910 = 10'h32e == io_inputs_0 ? 7'h64 : _GEN_4909; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4911 = 10'h32f == io_inputs_0 ? 7'h64 : _GEN_4910; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4912 = 10'h330 == io_inputs_0 ? 7'h64 : _GEN_4911; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4913 = 10'h331 == io_inputs_0 ? 7'h64 : _GEN_4912; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4914 = 10'h332 == io_inputs_0 ? 7'h64 : _GEN_4913; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4915 = 10'h333 == io_inputs_0 ? 7'h64 : _GEN_4914; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4916 = 10'h334 == io_inputs_0 ? 7'h64 : _GEN_4915; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4917 = 10'h335 == io_inputs_0 ? 7'h64 : _GEN_4916; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4918 = 10'h336 == io_inputs_0 ? 7'h64 : _GEN_4917; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4919 = 10'h337 == io_inputs_0 ? 7'h64 : _GEN_4918; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4920 = 10'h338 == io_inputs_0 ? 7'h64 : _GEN_4919; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4921 = 10'h339 == io_inputs_0 ? 7'h64 : _GEN_4920; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4922 = 10'h33a == io_inputs_0 ? 7'h64 : _GEN_4921; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4923 = 10'h33b == io_inputs_0 ? 7'h64 : _GEN_4922; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4924 = 10'h33c == io_inputs_0 ? 7'h64 : _GEN_4923; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4925 = 10'h33d == io_inputs_0 ? 7'h64 : _GEN_4924; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4926 = 10'h33e == io_inputs_0 ? 7'h64 : _GEN_4925; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4927 = 10'h33f == io_inputs_0 ? 7'h64 : _GEN_4926; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4928 = 10'h340 == io_inputs_0 ? 7'h64 : _GEN_4927; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4929 = 10'h341 == io_inputs_0 ? 7'h64 : _GEN_4928; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4930 = 10'h342 == io_inputs_0 ? 7'h64 : _GEN_4929; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4931 = 10'h343 == io_inputs_0 ? 7'h64 : _GEN_4930; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4932 = 10'h344 == io_inputs_0 ? 7'h64 : _GEN_4931; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4933 = 10'h345 == io_inputs_0 ? 7'h64 : _GEN_4932; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4934 = 10'h346 == io_inputs_0 ? 7'h64 : _GEN_4933; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4935 = 10'h347 == io_inputs_0 ? 7'h64 : _GEN_4934; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4936 = 10'h348 == io_inputs_0 ? 7'h64 : _GEN_4935; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4937 = 10'h349 == io_inputs_0 ? 7'h64 : _GEN_4936; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4938 = 10'h34a == io_inputs_0 ? 7'h64 : _GEN_4937; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4939 = 10'h34b == io_inputs_0 ? 7'h64 : _GEN_4938; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4940 = 10'h34c == io_inputs_0 ? 7'h64 : _GEN_4939; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4941 = 10'h34d == io_inputs_0 ? 7'h64 : _GEN_4940; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4942 = 10'h34e == io_inputs_0 ? 7'h64 : _GEN_4941; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4943 = 10'h34f == io_inputs_0 ? 7'h64 : _GEN_4942; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4944 = 10'h350 == io_inputs_0 ? 7'h64 : _GEN_4943; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4945 = 10'h351 == io_inputs_0 ? 7'h64 : _GEN_4944; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4946 = 10'h352 == io_inputs_0 ? 7'h64 : _GEN_4945; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4947 = 10'h353 == io_inputs_0 ? 7'h64 : _GEN_4946; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4948 = 10'h354 == io_inputs_0 ? 7'h64 : _GEN_4947; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4949 = 10'h355 == io_inputs_0 ? 7'h64 : _GEN_4948; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4950 = 10'h356 == io_inputs_0 ? 7'h64 : _GEN_4949; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4951 = 10'h357 == io_inputs_0 ? 7'h64 : _GEN_4950; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4952 = 10'h358 == io_inputs_0 ? 7'h64 : _GEN_4951; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4953 = 10'h359 == io_inputs_0 ? 7'h64 : _GEN_4952; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4954 = 10'h35a == io_inputs_0 ? 7'h64 : _GEN_4953; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4955 = 10'h35b == io_inputs_0 ? 7'h64 : _GEN_4954; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4956 = 10'h35c == io_inputs_0 ? 7'h64 : _GEN_4955; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4957 = 10'h35d == io_inputs_0 ? 7'h64 : _GEN_4956; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4958 = 10'h35e == io_inputs_0 ? 7'h64 : _GEN_4957; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4959 = 10'h35f == io_inputs_0 ? 7'h64 : _GEN_4958; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4960 = 10'h360 == io_inputs_0 ? 7'h64 : _GEN_4959; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4961 = 10'h361 == io_inputs_0 ? 7'h64 : _GEN_4960; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4962 = 10'h362 == io_inputs_0 ? 7'h64 : _GEN_4961; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4963 = 10'h363 == io_inputs_0 ? 7'h64 : _GEN_4962; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4964 = 10'h364 == io_inputs_0 ? 7'h64 : _GEN_4963; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4965 = 10'h365 == io_inputs_0 ? 7'h64 : _GEN_4964; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4966 = 10'h366 == io_inputs_0 ? 7'h64 : _GEN_4965; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4967 = 10'h367 == io_inputs_0 ? 7'h64 : _GEN_4966; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4968 = 10'h368 == io_inputs_0 ? 7'h64 : _GEN_4967; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4969 = 10'h369 == io_inputs_0 ? 7'h64 : _GEN_4968; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4970 = 10'h36a == io_inputs_0 ? 7'h64 : _GEN_4969; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4971 = 10'h36b == io_inputs_0 ? 7'h64 : _GEN_4970; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4972 = 10'h36c == io_inputs_0 ? 7'h64 : _GEN_4971; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4973 = 10'h36d == io_inputs_0 ? 7'h64 : _GEN_4972; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4974 = 10'h36e == io_inputs_0 ? 7'h64 : _GEN_4973; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4975 = 10'h36f == io_inputs_0 ? 7'h64 : _GEN_4974; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4976 = 10'h370 == io_inputs_0 ? 7'h64 : _GEN_4975; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4977 = 10'h371 == io_inputs_0 ? 7'h64 : _GEN_4976; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4978 = 10'h372 == io_inputs_0 ? 7'h64 : _GEN_4977; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4979 = 10'h373 == io_inputs_0 ? 7'h64 : _GEN_4978; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4980 = 10'h374 == io_inputs_0 ? 7'h64 : _GEN_4979; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4981 = 10'h375 == io_inputs_0 ? 7'h64 : _GEN_4980; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4982 = 10'h376 == io_inputs_0 ? 7'h64 : _GEN_4981; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4983 = 10'h377 == io_inputs_0 ? 7'h64 : _GEN_4982; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4984 = 10'h378 == io_inputs_0 ? 7'h64 : _GEN_4983; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4985 = 10'h379 == io_inputs_0 ? 7'h64 : _GEN_4984; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4986 = 10'h37a == io_inputs_0 ? 7'h64 : _GEN_4985; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4987 = 10'h37b == io_inputs_0 ? 7'h64 : _GEN_4986; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4988 = 10'h37c == io_inputs_0 ? 7'h64 : _GEN_4987; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4989 = 10'h37d == io_inputs_0 ? 7'h64 : _GEN_4988; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4990 = 10'h37e == io_inputs_0 ? 7'h64 : _GEN_4989; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4991 = 10'h37f == io_inputs_0 ? 7'h64 : _GEN_4990; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4992 = 10'h380 == io_inputs_0 ? 7'h64 : _GEN_4991; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4993 = 10'h381 == io_inputs_0 ? 7'h64 : _GEN_4992; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4994 = 10'h382 == io_inputs_0 ? 7'h64 : _GEN_4993; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4995 = 10'h383 == io_inputs_0 ? 7'h64 : _GEN_4994; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4996 = 10'h384 == io_inputs_0 ? 7'h64 : _GEN_4995; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4997 = 10'h385 == io_inputs_0 ? 7'h64 : _GEN_4996; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4998 = 10'h386 == io_inputs_0 ? 7'h64 : _GEN_4997; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_4999 = 10'h387 == io_inputs_0 ? 7'h64 : _GEN_4998; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5000 = 10'h388 == io_inputs_0 ? 7'h64 : _GEN_4999; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5001 = 10'h389 == io_inputs_0 ? 7'h64 : _GEN_5000; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5002 = 10'h38a == io_inputs_0 ? 7'h64 : _GEN_5001; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5003 = 10'h38b == io_inputs_0 ? 7'h64 : _GEN_5002; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5004 = 10'h38c == io_inputs_0 ? 7'h64 : _GEN_5003; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5005 = 10'h38d == io_inputs_0 ? 7'h64 : _GEN_5004; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5006 = 10'h38e == io_inputs_0 ? 7'h64 : _GEN_5005; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5007 = 10'h38f == io_inputs_0 ? 7'h64 : _GEN_5006; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5008 = 10'h390 == io_inputs_0 ? 7'h64 : _GEN_5007; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5009 = 10'h391 == io_inputs_0 ? 7'h64 : _GEN_5008; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5010 = 10'h392 == io_inputs_0 ? 7'h64 : _GEN_5009; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5011 = 10'h393 == io_inputs_0 ? 7'h64 : _GEN_5010; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5012 = 10'h394 == io_inputs_0 ? 7'h64 : _GEN_5011; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5013 = 10'h395 == io_inputs_0 ? 7'h64 : _GEN_5012; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5014 = 10'h396 == io_inputs_0 ? 7'h64 : _GEN_5013; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5015 = 10'h397 == io_inputs_0 ? 7'h64 : _GEN_5014; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5016 = 10'h398 == io_inputs_0 ? 7'h64 : _GEN_5015; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5017 = 10'h399 == io_inputs_0 ? 7'h64 : _GEN_5016; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5018 = 10'h39a == io_inputs_0 ? 7'h64 : _GEN_5017; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5019 = 10'h39b == io_inputs_0 ? 7'h64 : _GEN_5018; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5020 = 10'h39c == io_inputs_0 ? 7'h64 : _GEN_5019; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5021 = 10'h39d == io_inputs_0 ? 7'h64 : _GEN_5020; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5022 = 10'h39e == io_inputs_0 ? 7'h64 : _GEN_5021; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5023 = 10'h39f == io_inputs_0 ? 7'h64 : _GEN_5022; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5024 = 10'h3a0 == io_inputs_0 ? 7'h64 : _GEN_5023; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5025 = 10'h3a1 == io_inputs_0 ? 7'h64 : _GEN_5024; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5026 = 10'h3a2 == io_inputs_0 ? 7'h64 : _GEN_5025; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5027 = 10'h3a3 == io_inputs_0 ? 7'h64 : _GEN_5026; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5028 = 10'h3a4 == io_inputs_0 ? 7'h64 : _GEN_5027; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5029 = 10'h3a5 == io_inputs_0 ? 7'h64 : _GEN_5028; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5030 = 10'h3a6 == io_inputs_0 ? 7'h64 : _GEN_5029; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5031 = 10'h3a7 == io_inputs_0 ? 7'h64 : _GEN_5030; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5032 = 10'h3a8 == io_inputs_0 ? 7'h64 : _GEN_5031; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5033 = 10'h3a9 == io_inputs_0 ? 7'h64 : _GEN_5032; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5034 = 10'h3aa == io_inputs_0 ? 7'h64 : _GEN_5033; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5035 = 10'h3ab == io_inputs_0 ? 7'h64 : _GEN_5034; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5036 = 10'h3ac == io_inputs_0 ? 7'h64 : _GEN_5035; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5037 = 10'h3ad == io_inputs_0 ? 7'h64 : _GEN_5036; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5038 = 10'h3ae == io_inputs_0 ? 7'h64 : _GEN_5037; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5039 = 10'h3af == io_inputs_0 ? 7'h64 : _GEN_5038; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5040 = 10'h3b0 == io_inputs_0 ? 7'h64 : _GEN_5039; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5041 = 10'h3b1 == io_inputs_0 ? 7'h64 : _GEN_5040; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5042 = 10'h3b2 == io_inputs_0 ? 7'h64 : _GEN_5041; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5043 = 10'h3b3 == io_inputs_0 ? 7'h64 : _GEN_5042; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5044 = 10'h3b4 == io_inputs_0 ? 7'h64 : _GEN_5043; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5045 = 10'h3b5 == io_inputs_0 ? 7'h64 : _GEN_5044; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5046 = 10'h3b6 == io_inputs_0 ? 7'h64 : _GEN_5045; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5047 = 10'h3b7 == io_inputs_0 ? 7'h64 : _GEN_5046; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5048 = 10'h3b8 == io_inputs_0 ? 7'h64 : _GEN_5047; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5049 = 10'h3b9 == io_inputs_0 ? 7'h64 : _GEN_5048; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5050 = 10'h3ba == io_inputs_0 ? 7'h64 : _GEN_5049; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5051 = 10'h3bb == io_inputs_0 ? 7'h64 : _GEN_5050; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5052 = 10'h3bc == io_inputs_0 ? 7'h64 : _GEN_5051; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5053 = 10'h3bd == io_inputs_0 ? 7'h64 : _GEN_5052; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5054 = 10'h3be == io_inputs_0 ? 7'h64 : _GEN_5053; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5055 = 10'h3bf == io_inputs_0 ? 7'h64 : _GEN_5054; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5056 = 10'h3c0 == io_inputs_0 ? 7'h64 : _GEN_5055; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5057 = 10'h3c1 == io_inputs_0 ? 7'h64 : _GEN_5056; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5058 = 10'h3c2 == io_inputs_0 ? 7'h64 : _GEN_5057; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5059 = 10'h3c3 == io_inputs_0 ? 7'h64 : _GEN_5058; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5060 = 10'h3c4 == io_inputs_0 ? 7'h64 : _GEN_5059; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5061 = 10'h3c5 == io_inputs_0 ? 7'h64 : _GEN_5060; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5062 = 10'h3c6 == io_inputs_0 ? 7'h64 : _GEN_5061; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5063 = 10'h3c7 == io_inputs_0 ? 7'h64 : _GEN_5062; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5064 = 10'h3c8 == io_inputs_0 ? 7'h64 : _GEN_5063; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5065 = 10'h3c9 == io_inputs_0 ? 7'h64 : _GEN_5064; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5066 = 10'h3ca == io_inputs_0 ? 7'h64 : _GEN_5065; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5067 = 10'h3cb == io_inputs_0 ? 7'h64 : _GEN_5066; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5068 = 10'h3cc == io_inputs_0 ? 7'h64 : _GEN_5067; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5069 = 10'h3cd == io_inputs_0 ? 7'h64 : _GEN_5068; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5070 = 10'h3ce == io_inputs_0 ? 7'h64 : _GEN_5069; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5071 = 10'h3cf == io_inputs_0 ? 7'h64 : _GEN_5070; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5072 = 10'h3d0 == io_inputs_0 ? 7'h64 : _GEN_5071; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5073 = 10'h3d1 == io_inputs_0 ? 7'h64 : _GEN_5072; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5074 = 10'h3d2 == io_inputs_0 ? 7'h64 : _GEN_5073; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5075 = 10'h3d3 == io_inputs_0 ? 7'h64 : _GEN_5074; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5076 = 10'h3d4 == io_inputs_0 ? 7'h64 : _GEN_5075; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5077 = 10'h3d5 == io_inputs_0 ? 7'h64 : _GEN_5076; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5078 = 10'h3d6 == io_inputs_0 ? 7'h64 : _GEN_5077; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5079 = 10'h3d7 == io_inputs_0 ? 7'h64 : _GEN_5078; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5080 = 10'h3d8 == io_inputs_0 ? 7'h64 : _GEN_5079; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5081 = 10'h3d9 == io_inputs_0 ? 7'h64 : _GEN_5080; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5082 = 10'h3da == io_inputs_0 ? 7'h64 : _GEN_5081; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5083 = 10'h3db == io_inputs_0 ? 7'h64 : _GEN_5082; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5084 = 10'h3dc == io_inputs_0 ? 7'h64 : _GEN_5083; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5085 = 10'h3dd == io_inputs_0 ? 7'h64 : _GEN_5084; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5086 = 10'h3de == io_inputs_0 ? 7'h64 : _GEN_5085; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5087 = 10'h3df == io_inputs_0 ? 7'h64 : _GEN_5086; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5088 = 10'h3e0 == io_inputs_0 ? 7'h64 : _GEN_5087; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5089 = 10'h3e1 == io_inputs_0 ? 7'h64 : _GEN_5088; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5090 = 10'h3e2 == io_inputs_0 ? 7'h64 : _GEN_5089; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5091 = 10'h3e3 == io_inputs_0 ? 7'h64 : _GEN_5090; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5092 = 10'h3e4 == io_inputs_0 ? 7'h64 : _GEN_5091; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5093 = 10'h3e5 == io_inputs_0 ? 7'h64 : _GEN_5092; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5094 = 10'h3e6 == io_inputs_0 ? 7'h64 : _GEN_5093; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5095 = 10'h3e7 == io_inputs_0 ? 7'h64 : _GEN_5094; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5096 = 10'h3e8 == io_inputs_0 ? 7'h64 : _GEN_5095; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5097 = 10'h3e9 == io_inputs_0 ? 7'h64 : _GEN_5096; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5098 = 10'h3ea == io_inputs_0 ? 7'h64 : _GEN_5097; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5099 = 10'h3eb == io_inputs_0 ? 7'h64 : _GEN_5098; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5100 = 10'h3ec == io_inputs_0 ? 7'h64 : _GEN_5099; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5101 = 10'h3ed == io_inputs_0 ? 7'h64 : _GEN_5100; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5102 = 10'h3ee == io_inputs_0 ? 7'h64 : _GEN_5101; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5103 = 10'h3ef == io_inputs_0 ? 7'h64 : _GEN_5102; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5104 = 10'h3f0 == io_inputs_0 ? 7'h64 : _GEN_5103; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5105 = 10'h3f1 == io_inputs_0 ? 7'h64 : _GEN_5104; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5106 = 10'h3f2 == io_inputs_0 ? 7'h64 : _GEN_5105; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5107 = 10'h3f3 == io_inputs_0 ? 7'h64 : _GEN_5106; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5108 = 10'h3f4 == io_inputs_0 ? 7'h64 : _GEN_5107; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5109 = 10'h3f5 == io_inputs_0 ? 7'h64 : _GEN_5108; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5110 = 10'h3f6 == io_inputs_0 ? 7'h64 : _GEN_5109; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5111 = 10'h3f7 == io_inputs_0 ? 7'h64 : _GEN_5110; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5112 = 10'h3f8 == io_inputs_0 ? 7'h64 : _GEN_5111; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5113 = 10'h3f9 == io_inputs_0 ? 7'h64 : _GEN_5112; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5114 = 10'h3fa == io_inputs_0 ? 7'h64 : _GEN_5113; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5115 = 10'h3fb == io_inputs_0 ? 7'h64 : _GEN_5114; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5116 = 10'h3fc == io_inputs_0 ? 7'h64 : _GEN_5115; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5141 = 8'h15 == io_inputs_1[7:0] ? 7'h5f : 7'h64; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5142 = 8'h16 == io_inputs_1[7:0] ? 7'h5a : _GEN_5141; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5143 = 8'h17 == io_inputs_1[7:0] ? 7'h55 : _GEN_5142; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5144 = 8'h18 == io_inputs_1[7:0] ? 7'h50 : _GEN_5143; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5145 = 8'h19 == io_inputs_1[7:0] ? 7'h4b : _GEN_5144; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5146 = 8'h1a == io_inputs_1[7:0] ? 7'h46 : _GEN_5145; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5147 = 8'h1b == io_inputs_1[7:0] ? 7'h41 : _GEN_5146; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5148 = 8'h1c == io_inputs_1[7:0] ? 7'h3c : _GEN_5147; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5149 = 8'h1d == io_inputs_1[7:0] ? 7'h37 : _GEN_5148; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5150 = 8'h1e == io_inputs_1[7:0] ? 7'h32 : _GEN_5149; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5151 = 8'h1f == io_inputs_1[7:0] ? 7'h2d : _GEN_5150; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5152 = 8'h20 == io_inputs_1[7:0] ? 7'h28 : _GEN_5151; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5153 = 8'h21 == io_inputs_1[7:0] ? 7'h23 : _GEN_5152; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5154 = 8'h22 == io_inputs_1[7:0] ? 7'h1e : _GEN_5153; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5155 = 8'h23 == io_inputs_1[7:0] ? 7'h19 : _GEN_5154; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5156 = 8'h24 == io_inputs_1[7:0] ? 7'h14 : _GEN_5155; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5157 = 8'h25 == io_inputs_1[7:0] ? 7'hf : _GEN_5156; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5158 = 8'h26 == io_inputs_1[7:0] ? 7'ha : _GEN_5157; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5159 = 8'h27 == io_inputs_1[7:0] ? 7'h5 : _GEN_5158; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5160 = 8'h28 == io_inputs_1[7:0] ? 7'h0 : _GEN_5159; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5161 = 8'h29 == io_inputs_1[7:0] ? 7'h0 : _GEN_5160; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5162 = 8'h2a == io_inputs_1[7:0] ? 7'h0 : _GEN_5161; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5163 = 8'h2b == io_inputs_1[7:0] ? 7'h0 : _GEN_5162; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5164 = 8'h2c == io_inputs_1[7:0] ? 7'h0 : _GEN_5163; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5165 = 8'h2d == io_inputs_1[7:0] ? 7'h0 : _GEN_5164; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5166 = 8'h2e == io_inputs_1[7:0] ? 7'h0 : _GEN_5165; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5167 = 8'h2f == io_inputs_1[7:0] ? 7'h0 : _GEN_5166; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5168 = 8'h30 == io_inputs_1[7:0] ? 7'h0 : _GEN_5167; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5169 = 8'h31 == io_inputs_1[7:0] ? 7'h0 : _GEN_5168; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5170 = 8'h32 == io_inputs_1[7:0] ? 7'h0 : _GEN_5169; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5171 = 8'h33 == io_inputs_1[7:0] ? 7'h0 : _GEN_5170; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5172 = 8'h34 == io_inputs_1[7:0] ? 7'h0 : _GEN_5171; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5173 = 8'h35 == io_inputs_1[7:0] ? 7'h0 : _GEN_5172; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5174 = 8'h36 == io_inputs_1[7:0] ? 7'h0 : _GEN_5173; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5175 = 8'h37 == io_inputs_1[7:0] ? 7'h0 : _GEN_5174; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5176 = 8'h38 == io_inputs_1[7:0] ? 7'h0 : _GEN_5175; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5177 = 8'h39 == io_inputs_1[7:0] ? 7'h0 : _GEN_5176; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5178 = 8'h3a == io_inputs_1[7:0] ? 7'h0 : _GEN_5177; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5179 = 8'h3b == io_inputs_1[7:0] ? 7'h0 : _GEN_5178; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5180 = 8'h3c == io_inputs_1[7:0] ? 7'h0 : _GEN_5179; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5181 = 8'h3d == io_inputs_1[7:0] ? 7'h0 : _GEN_5180; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5182 = 8'h3e == io_inputs_1[7:0] ? 7'h0 : _GEN_5181; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5183 = 8'h3f == io_inputs_1[7:0] ? 7'h0 : _GEN_5182; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5184 = 8'h40 == io_inputs_1[7:0] ? 7'h0 : _GEN_5183; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5185 = 8'h41 == io_inputs_1[7:0] ? 7'h0 : _GEN_5184; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5186 = 8'h42 == io_inputs_1[7:0] ? 7'h0 : _GEN_5185; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5187 = 8'h43 == io_inputs_1[7:0] ? 7'h0 : _GEN_5186; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5188 = 8'h44 == io_inputs_1[7:0] ? 7'h0 : _GEN_5187; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5189 = 8'h45 == io_inputs_1[7:0] ? 7'h0 : _GEN_5188; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5190 = 8'h46 == io_inputs_1[7:0] ? 7'h0 : _GEN_5189; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5191 = 8'h47 == io_inputs_1[7:0] ? 7'h0 : _GEN_5190; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5192 = 8'h48 == io_inputs_1[7:0] ? 7'h0 : _GEN_5191; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5193 = 8'h49 == io_inputs_1[7:0] ? 7'h0 : _GEN_5192; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5194 = 8'h4a == io_inputs_1[7:0] ? 7'h0 : _GEN_5193; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5195 = 8'h4b == io_inputs_1[7:0] ? 7'h0 : _GEN_5194; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5196 = 8'h4c == io_inputs_1[7:0] ? 7'h0 : _GEN_5195; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5197 = 8'h4d == io_inputs_1[7:0] ? 7'h0 : _GEN_5196; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5198 = 8'h4e == io_inputs_1[7:0] ? 7'h0 : _GEN_5197; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5199 = 8'h4f == io_inputs_1[7:0] ? 7'h0 : _GEN_5198; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5200 = 8'h50 == io_inputs_1[7:0] ? 7'h0 : _GEN_5199; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5201 = 8'h51 == io_inputs_1[7:0] ? 7'h0 : _GEN_5200; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5202 = 8'h52 == io_inputs_1[7:0] ? 7'h0 : _GEN_5201; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5203 = 8'h53 == io_inputs_1[7:0] ? 7'h0 : _GEN_5202; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5204 = 8'h54 == io_inputs_1[7:0] ? 7'h0 : _GEN_5203; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5205 = 8'h55 == io_inputs_1[7:0] ? 7'h0 : _GEN_5204; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5206 = 8'h56 == io_inputs_1[7:0] ? 7'h0 : _GEN_5205; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5207 = 8'h57 == io_inputs_1[7:0] ? 7'h0 : _GEN_5206; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5208 = 8'h58 == io_inputs_1[7:0] ? 7'h0 : _GEN_5207; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5209 = 8'h59 == io_inputs_1[7:0] ? 7'h0 : _GEN_5208; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5210 = 8'h5a == io_inputs_1[7:0] ? 7'h0 : _GEN_5209; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5211 = 8'h5b == io_inputs_1[7:0] ? 7'h0 : _GEN_5210; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5212 = 8'h5c == io_inputs_1[7:0] ? 7'h0 : _GEN_5211; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5213 = 8'h5d == io_inputs_1[7:0] ? 7'h0 : _GEN_5212; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5214 = 8'h5e == io_inputs_1[7:0] ? 7'h0 : _GEN_5213; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5215 = 8'h5f == io_inputs_1[7:0] ? 7'h0 : _GEN_5214; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5216 = 8'h60 == io_inputs_1[7:0] ? 7'h0 : _GEN_5215; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5217 = 8'h61 == io_inputs_1[7:0] ? 7'h0 : _GEN_5216; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5218 = 8'h62 == io_inputs_1[7:0] ? 7'h0 : _GEN_5217; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5219 = 8'h63 == io_inputs_1[7:0] ? 7'h0 : _GEN_5218; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5220 = 8'h64 == io_inputs_1[7:0] ? 7'h0 : _GEN_5219; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5221 = 8'h65 == io_inputs_1[7:0] ? 7'h0 : _GEN_5220; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5222 = 8'h66 == io_inputs_1[7:0] ? 7'h0 : _GEN_5221; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5223 = 8'h67 == io_inputs_1[7:0] ? 7'h0 : _GEN_5222; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5224 = 8'h68 == io_inputs_1[7:0] ? 7'h0 : _GEN_5223; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5225 = 8'h69 == io_inputs_1[7:0] ? 7'h0 : _GEN_5224; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5226 = 8'h6a == io_inputs_1[7:0] ? 7'h0 : _GEN_5225; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5227 = 8'h6b == io_inputs_1[7:0] ? 7'h0 : _GEN_5226; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5228 = 8'h6c == io_inputs_1[7:0] ? 7'h0 : _GEN_5227; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5229 = 8'h6d == io_inputs_1[7:0] ? 7'h0 : _GEN_5228; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5230 = 8'h6e == io_inputs_1[7:0] ? 7'h0 : _GEN_5229; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5231 = 8'h6f == io_inputs_1[7:0] ? 7'h0 : _GEN_5230; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5232 = 8'h70 == io_inputs_1[7:0] ? 7'h0 : _GEN_5231; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5233 = 8'h71 == io_inputs_1[7:0] ? 7'h0 : _GEN_5232; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5234 = 8'h72 == io_inputs_1[7:0] ? 7'h0 : _GEN_5233; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5235 = 8'h73 == io_inputs_1[7:0] ? 7'h0 : _GEN_5234; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5236 = 8'h74 == io_inputs_1[7:0] ? 7'h0 : _GEN_5235; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5237 = 8'h75 == io_inputs_1[7:0] ? 7'h0 : _GEN_5236; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5238 = 8'h76 == io_inputs_1[7:0] ? 7'h0 : _GEN_5237; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5239 = 8'h77 == io_inputs_1[7:0] ? 7'h0 : _GEN_5238; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5240 = 8'h78 == io_inputs_1[7:0] ? 7'h0 : _GEN_5239; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5241 = 8'h79 == io_inputs_1[7:0] ? 7'h0 : _GEN_5240; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5242 = 8'h7a == io_inputs_1[7:0] ? 7'h0 : _GEN_5241; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5243 = 8'h7b == io_inputs_1[7:0] ? 7'h0 : _GEN_5242; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5244 = 8'h7c == io_inputs_1[7:0] ? 7'h0 : _GEN_5243; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5245 = 8'h7d == io_inputs_1[7:0] ? 7'h0 : _GEN_5244; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5246 = 8'h7e == io_inputs_1[7:0] ? 7'h0 : _GEN_5245; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5247 = 8'h7f == io_inputs_1[7:0] ? 7'h0 : _GEN_5246; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5248 = 8'h80 == io_inputs_1[7:0] ? 7'h0 : _GEN_5247; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5249 = 8'h81 == io_inputs_1[7:0] ? 7'h0 : _GEN_5248; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5250 = 8'h82 == io_inputs_1[7:0] ? 7'h0 : _GEN_5249; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5251 = 8'h83 == io_inputs_1[7:0] ? 7'h0 : _GEN_5250; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5252 = 8'h84 == io_inputs_1[7:0] ? 7'h0 : _GEN_5251; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5253 = 8'h85 == io_inputs_1[7:0] ? 7'h0 : _GEN_5252; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5254 = 8'h86 == io_inputs_1[7:0] ? 7'h0 : _GEN_5253; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5255 = 8'h87 == io_inputs_1[7:0] ? 7'h0 : _GEN_5254; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5256 = 8'h88 == io_inputs_1[7:0] ? 7'h0 : _GEN_5255; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5257 = 8'h89 == io_inputs_1[7:0] ? 7'h0 : _GEN_5256; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5258 = 8'h8a == io_inputs_1[7:0] ? 7'h0 : _GEN_5257; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5259 = 8'h8b == io_inputs_1[7:0] ? 7'h0 : _GEN_5258; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5260 = 8'h8c == io_inputs_1[7:0] ? 7'h0 : _GEN_5259; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5261 = 8'h8d == io_inputs_1[7:0] ? 7'h0 : _GEN_5260; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5262 = 8'h8e == io_inputs_1[7:0] ? 7'h0 : _GEN_5261; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5263 = 8'h8f == io_inputs_1[7:0] ? 7'h0 : _GEN_5262; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5264 = 8'h90 == io_inputs_1[7:0] ? 7'h0 : _GEN_5263; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5265 = 8'h91 == io_inputs_1[7:0] ? 7'h0 : _GEN_5264; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5266 = 8'h92 == io_inputs_1[7:0] ? 7'h0 : _GEN_5265; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5267 = 8'h93 == io_inputs_1[7:0] ? 7'h0 : _GEN_5266; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5268 = 8'h94 == io_inputs_1[7:0] ? 7'h0 : _GEN_5267; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5269 = 8'h95 == io_inputs_1[7:0] ? 7'h0 : _GEN_5268; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5270 = 8'h96 == io_inputs_1[7:0] ? 7'h0 : _GEN_5269; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5271 = 8'h97 == io_inputs_1[7:0] ? 7'h0 : _GEN_5270; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5272 = 8'h98 == io_inputs_1[7:0] ? 7'h0 : _GEN_5271; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5273 = 8'h99 == io_inputs_1[7:0] ? 7'h0 : _GEN_5272; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5274 = 8'h9a == io_inputs_1[7:0] ? 7'h0 : _GEN_5273; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5275 = 8'h9b == io_inputs_1[7:0] ? 7'h0 : _GEN_5274; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5276 = 8'h9c == io_inputs_1[7:0] ? 7'h0 : _GEN_5275; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5277 = 8'h9d == io_inputs_1[7:0] ? 7'h0 : _GEN_5276; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5278 = 8'h9e == io_inputs_1[7:0] ? 7'h0 : _GEN_5277; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5279 = 8'h9f == io_inputs_1[7:0] ? 7'h0 : _GEN_5278; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5280 = 8'ha0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5279; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5281 = 8'ha1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5280; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5282 = 8'ha2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5281; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5283 = 8'ha3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5282; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5284 = 8'ha4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5283; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5285 = 8'ha5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5284; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5286 = 8'ha6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5285; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5287 = 8'ha7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5286; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5288 = 8'ha8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5287; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5289 = 8'ha9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5288; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5290 = 8'haa == io_inputs_1[7:0] ? 7'h0 : _GEN_5289; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5291 = 8'hab == io_inputs_1[7:0] ? 7'h0 : _GEN_5290; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5292 = 8'hac == io_inputs_1[7:0] ? 7'h0 : _GEN_5291; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5293 = 8'had == io_inputs_1[7:0] ? 7'h0 : _GEN_5292; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5294 = 8'hae == io_inputs_1[7:0] ? 7'h0 : _GEN_5293; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5295 = 8'haf == io_inputs_1[7:0] ? 7'h0 : _GEN_5294; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5296 = 8'hb0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5295; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5297 = 8'hb1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5296; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5298 = 8'hb2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5297; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5299 = 8'hb3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5298; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5300 = 8'hb4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5299; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5301 = 8'hb5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5300; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5302 = 8'hb6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5301; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5303 = 8'hb7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5302; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5304 = 8'hb8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5303; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5305 = 8'hb9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5304; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5306 = 8'hba == io_inputs_1[7:0] ? 7'h0 : _GEN_5305; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5307 = 8'hbb == io_inputs_1[7:0] ? 7'h0 : _GEN_5306; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5308 = 8'hbc == io_inputs_1[7:0] ? 7'h0 : _GEN_5307; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5309 = 8'hbd == io_inputs_1[7:0] ? 7'h0 : _GEN_5308; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5310 = 8'hbe == io_inputs_1[7:0] ? 7'h0 : _GEN_5309; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5311 = 8'hbf == io_inputs_1[7:0] ? 7'h0 : _GEN_5310; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5312 = 8'hc0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5311; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5313 = 8'hc1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5312; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5314 = 8'hc2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5313; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5315 = 8'hc3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5314; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5316 = 8'hc4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5315; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5317 = 8'hc5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5316; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5318 = 8'hc6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5317; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5319 = 8'hc7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5318; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5320 = 8'hc8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5319; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5321 = 8'hc9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5320; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5322 = 8'hca == io_inputs_1[7:0] ? 7'h0 : _GEN_5321; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5323 = 8'hcb == io_inputs_1[7:0] ? 7'h0 : _GEN_5322; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5324 = 8'hcc == io_inputs_1[7:0] ? 7'h0 : _GEN_5323; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5325 = 8'hcd == io_inputs_1[7:0] ? 7'h0 : _GEN_5324; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5326 = 8'hce == io_inputs_1[7:0] ? 7'h0 : _GEN_5325; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5327 = 8'hcf == io_inputs_1[7:0] ? 7'h0 : _GEN_5326; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5328 = 8'hd0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5327; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5329 = 8'hd1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5328; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5330 = 8'hd2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5329; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5331 = 8'hd3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5330; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5332 = 8'hd4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5331; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5333 = 8'hd5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5332; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5334 = 8'hd6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5333; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5335 = 8'hd7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5334; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5336 = 8'hd8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5335; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5337 = 8'hd9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5336; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5338 = 8'hda == io_inputs_1[7:0] ? 7'h0 : _GEN_5337; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5339 = 8'hdb == io_inputs_1[7:0] ? 7'h0 : _GEN_5338; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5340 = 8'hdc == io_inputs_1[7:0] ? 7'h0 : _GEN_5339; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5341 = 8'hdd == io_inputs_1[7:0] ? 7'h0 : _GEN_5340; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5342 = 8'hde == io_inputs_1[7:0] ? 7'h0 : _GEN_5341; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5343 = 8'hdf == io_inputs_1[7:0] ? 7'h0 : _GEN_5342; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5344 = 8'he0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5343; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5345 = 8'he1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5344; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5346 = 8'he2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5345; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5347 = 8'he3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5346; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5348 = 8'he4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5347; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5349 = 8'he5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5348; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5350 = 8'he6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5349; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5351 = 8'he7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5350; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5352 = 8'he8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5351; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5353 = 8'he9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5352; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5354 = 8'hea == io_inputs_1[7:0] ? 7'h0 : _GEN_5353; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5355 = 8'heb == io_inputs_1[7:0] ? 7'h0 : _GEN_5354; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5356 = 8'hec == io_inputs_1[7:0] ? 7'h0 : _GEN_5355; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5357 = 8'hed == io_inputs_1[7:0] ? 7'h0 : _GEN_5356; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5358 = 8'hee == io_inputs_1[7:0] ? 7'h0 : _GEN_5357; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5359 = 8'hef == io_inputs_1[7:0] ? 7'h0 : _GEN_5358; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5360 = 8'hf0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5359; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5361 = 8'hf1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5360; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5362 = 8'hf2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5361; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5363 = 8'hf3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5362; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5364 = 8'hf4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5363; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5365 = 8'hf5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5364; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5366 = 8'hf6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5365; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5367 = 8'hf7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5366; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5368 = 8'hf8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5367; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5369 = 8'hf9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5368; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5370 = 8'hfa == io_inputs_1[7:0] ? 7'h0 : _GEN_5369; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5371 = 8'hfb == io_inputs_1[7:0] ? 7'h0 : _GEN_5370; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5372 = 8'hfc == io_inputs_1[7:0] ? 7'h0 : _GEN_5371; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5397 = 8'h15 == io_inputs_1[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5398 = 8'h16 == io_inputs_1[7:0] ? 7'ha : _GEN_5397; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5399 = 8'h17 == io_inputs_1[7:0] ? 7'hf : _GEN_5398; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5400 = 8'h18 == io_inputs_1[7:0] ? 7'h14 : _GEN_5399; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5401 = 8'h19 == io_inputs_1[7:0] ? 7'h19 : _GEN_5400; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5402 = 8'h1a == io_inputs_1[7:0] ? 7'h1e : _GEN_5401; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5403 = 8'h1b == io_inputs_1[7:0] ? 7'h23 : _GEN_5402; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5404 = 8'h1c == io_inputs_1[7:0] ? 7'h28 : _GEN_5403; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5405 = 8'h1d == io_inputs_1[7:0] ? 7'h2d : _GEN_5404; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5406 = 8'h1e == io_inputs_1[7:0] ? 7'h32 : _GEN_5405; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5407 = 8'h1f == io_inputs_1[7:0] ? 7'h37 : _GEN_5406; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5408 = 8'h20 == io_inputs_1[7:0] ? 7'h3c : _GEN_5407; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5409 = 8'h21 == io_inputs_1[7:0] ? 7'h41 : _GEN_5408; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5410 = 8'h22 == io_inputs_1[7:0] ? 7'h46 : _GEN_5409; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5411 = 8'h23 == io_inputs_1[7:0] ? 7'h4b : _GEN_5410; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5412 = 8'h24 == io_inputs_1[7:0] ? 7'h50 : _GEN_5411; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5413 = 8'h25 == io_inputs_1[7:0] ? 7'h55 : _GEN_5412; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5414 = 8'h26 == io_inputs_1[7:0] ? 7'h5a : _GEN_5413; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5415 = 8'h27 == io_inputs_1[7:0] ? 7'h5f : _GEN_5414; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5416 = 8'h28 == io_inputs_1[7:0] ? 7'h64 : _GEN_5415; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5417 = 8'h29 == io_inputs_1[7:0] ? 7'h64 : _GEN_5416; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5418 = 8'h2a == io_inputs_1[7:0] ? 7'h64 : _GEN_5417; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5419 = 8'h2b == io_inputs_1[7:0] ? 7'h64 : _GEN_5418; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5420 = 8'h2c == io_inputs_1[7:0] ? 7'h64 : _GEN_5419; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5421 = 8'h2d == io_inputs_1[7:0] ? 7'h64 : _GEN_5420; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5422 = 8'h2e == io_inputs_1[7:0] ? 7'h64 : _GEN_5421; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5423 = 8'h2f == io_inputs_1[7:0] ? 7'h64 : _GEN_5422; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5424 = 8'h30 == io_inputs_1[7:0] ? 7'h64 : _GEN_5423; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5425 = 8'h31 == io_inputs_1[7:0] ? 7'h64 : _GEN_5424; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5426 = 8'h32 == io_inputs_1[7:0] ? 7'h64 : _GEN_5425; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5427 = 8'h33 == io_inputs_1[7:0] ? 7'h64 : _GEN_5426; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5428 = 8'h34 == io_inputs_1[7:0] ? 7'h64 : _GEN_5427; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5429 = 8'h35 == io_inputs_1[7:0] ? 7'h64 : _GEN_5428; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5430 = 8'h36 == io_inputs_1[7:0] ? 7'h64 : _GEN_5429; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5431 = 8'h37 == io_inputs_1[7:0] ? 7'h64 : _GEN_5430; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5432 = 8'h38 == io_inputs_1[7:0] ? 7'h64 : _GEN_5431; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5433 = 8'h39 == io_inputs_1[7:0] ? 7'h64 : _GEN_5432; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5434 = 8'h3a == io_inputs_1[7:0] ? 7'h64 : _GEN_5433; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5435 = 8'h3b == io_inputs_1[7:0] ? 7'h64 : _GEN_5434; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5436 = 8'h3c == io_inputs_1[7:0] ? 7'h64 : _GEN_5435; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5437 = 8'h3d == io_inputs_1[7:0] ? 7'h5f : _GEN_5436; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5438 = 8'h3e == io_inputs_1[7:0] ? 7'h5a : _GEN_5437; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5439 = 8'h3f == io_inputs_1[7:0] ? 7'h55 : _GEN_5438; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5440 = 8'h40 == io_inputs_1[7:0] ? 7'h50 : _GEN_5439; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5441 = 8'h41 == io_inputs_1[7:0] ? 7'h4b : _GEN_5440; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5442 = 8'h42 == io_inputs_1[7:0] ? 7'h46 : _GEN_5441; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5443 = 8'h43 == io_inputs_1[7:0] ? 7'h41 : _GEN_5442; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5444 = 8'h44 == io_inputs_1[7:0] ? 7'h3c : _GEN_5443; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5445 = 8'h45 == io_inputs_1[7:0] ? 7'h37 : _GEN_5444; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5446 = 8'h46 == io_inputs_1[7:0] ? 7'h32 : _GEN_5445; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5447 = 8'h47 == io_inputs_1[7:0] ? 7'h2d : _GEN_5446; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5448 = 8'h48 == io_inputs_1[7:0] ? 7'h28 : _GEN_5447; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5449 = 8'h49 == io_inputs_1[7:0] ? 7'h23 : _GEN_5448; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5450 = 8'h4a == io_inputs_1[7:0] ? 7'h1e : _GEN_5449; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5451 = 8'h4b == io_inputs_1[7:0] ? 7'h19 : _GEN_5450; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5452 = 8'h4c == io_inputs_1[7:0] ? 7'h14 : _GEN_5451; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5453 = 8'h4d == io_inputs_1[7:0] ? 7'hf : _GEN_5452; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5454 = 8'h4e == io_inputs_1[7:0] ? 7'ha : _GEN_5453; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5455 = 8'h4f == io_inputs_1[7:0] ? 7'h5 : _GEN_5454; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5456 = 8'h50 == io_inputs_1[7:0] ? 7'h0 : _GEN_5455; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5457 = 8'h51 == io_inputs_1[7:0] ? 7'h0 : _GEN_5456; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5458 = 8'h52 == io_inputs_1[7:0] ? 7'h0 : _GEN_5457; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5459 = 8'h53 == io_inputs_1[7:0] ? 7'h0 : _GEN_5458; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5460 = 8'h54 == io_inputs_1[7:0] ? 7'h0 : _GEN_5459; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5461 = 8'h55 == io_inputs_1[7:0] ? 7'h0 : _GEN_5460; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5462 = 8'h56 == io_inputs_1[7:0] ? 7'h0 : _GEN_5461; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5463 = 8'h57 == io_inputs_1[7:0] ? 7'h0 : _GEN_5462; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5464 = 8'h58 == io_inputs_1[7:0] ? 7'h0 : _GEN_5463; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5465 = 8'h59 == io_inputs_1[7:0] ? 7'h0 : _GEN_5464; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5466 = 8'h5a == io_inputs_1[7:0] ? 7'h0 : _GEN_5465; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5467 = 8'h5b == io_inputs_1[7:0] ? 7'h0 : _GEN_5466; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5468 = 8'h5c == io_inputs_1[7:0] ? 7'h0 : _GEN_5467; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5469 = 8'h5d == io_inputs_1[7:0] ? 7'h0 : _GEN_5468; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5470 = 8'h5e == io_inputs_1[7:0] ? 7'h0 : _GEN_5469; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5471 = 8'h5f == io_inputs_1[7:0] ? 7'h0 : _GEN_5470; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5472 = 8'h60 == io_inputs_1[7:0] ? 7'h0 : _GEN_5471; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5473 = 8'h61 == io_inputs_1[7:0] ? 7'h0 : _GEN_5472; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5474 = 8'h62 == io_inputs_1[7:0] ? 7'h0 : _GEN_5473; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5475 = 8'h63 == io_inputs_1[7:0] ? 7'h0 : _GEN_5474; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5476 = 8'h64 == io_inputs_1[7:0] ? 7'h0 : _GEN_5475; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5477 = 8'h65 == io_inputs_1[7:0] ? 7'h0 : _GEN_5476; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5478 = 8'h66 == io_inputs_1[7:0] ? 7'h0 : _GEN_5477; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5479 = 8'h67 == io_inputs_1[7:0] ? 7'h0 : _GEN_5478; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5480 = 8'h68 == io_inputs_1[7:0] ? 7'h0 : _GEN_5479; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5481 = 8'h69 == io_inputs_1[7:0] ? 7'h0 : _GEN_5480; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5482 = 8'h6a == io_inputs_1[7:0] ? 7'h0 : _GEN_5481; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5483 = 8'h6b == io_inputs_1[7:0] ? 7'h0 : _GEN_5482; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5484 = 8'h6c == io_inputs_1[7:0] ? 7'h0 : _GEN_5483; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5485 = 8'h6d == io_inputs_1[7:0] ? 7'h0 : _GEN_5484; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5486 = 8'h6e == io_inputs_1[7:0] ? 7'h0 : _GEN_5485; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5487 = 8'h6f == io_inputs_1[7:0] ? 7'h0 : _GEN_5486; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5488 = 8'h70 == io_inputs_1[7:0] ? 7'h0 : _GEN_5487; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5489 = 8'h71 == io_inputs_1[7:0] ? 7'h0 : _GEN_5488; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5490 = 8'h72 == io_inputs_1[7:0] ? 7'h0 : _GEN_5489; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5491 = 8'h73 == io_inputs_1[7:0] ? 7'h0 : _GEN_5490; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5492 = 8'h74 == io_inputs_1[7:0] ? 7'h0 : _GEN_5491; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5493 = 8'h75 == io_inputs_1[7:0] ? 7'h0 : _GEN_5492; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5494 = 8'h76 == io_inputs_1[7:0] ? 7'h0 : _GEN_5493; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5495 = 8'h77 == io_inputs_1[7:0] ? 7'h0 : _GEN_5494; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5496 = 8'h78 == io_inputs_1[7:0] ? 7'h0 : _GEN_5495; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5497 = 8'h79 == io_inputs_1[7:0] ? 7'h0 : _GEN_5496; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5498 = 8'h7a == io_inputs_1[7:0] ? 7'h0 : _GEN_5497; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5499 = 8'h7b == io_inputs_1[7:0] ? 7'h0 : _GEN_5498; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5500 = 8'h7c == io_inputs_1[7:0] ? 7'h0 : _GEN_5499; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5501 = 8'h7d == io_inputs_1[7:0] ? 7'h0 : _GEN_5500; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5502 = 8'h7e == io_inputs_1[7:0] ? 7'h0 : _GEN_5501; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5503 = 8'h7f == io_inputs_1[7:0] ? 7'h0 : _GEN_5502; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5504 = 8'h80 == io_inputs_1[7:0] ? 7'h0 : _GEN_5503; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5505 = 8'h81 == io_inputs_1[7:0] ? 7'h0 : _GEN_5504; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5506 = 8'h82 == io_inputs_1[7:0] ? 7'h0 : _GEN_5505; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5507 = 8'h83 == io_inputs_1[7:0] ? 7'h0 : _GEN_5506; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5508 = 8'h84 == io_inputs_1[7:0] ? 7'h0 : _GEN_5507; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5509 = 8'h85 == io_inputs_1[7:0] ? 7'h0 : _GEN_5508; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5510 = 8'h86 == io_inputs_1[7:0] ? 7'h0 : _GEN_5509; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5511 = 8'h87 == io_inputs_1[7:0] ? 7'h0 : _GEN_5510; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5512 = 8'h88 == io_inputs_1[7:0] ? 7'h0 : _GEN_5511; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5513 = 8'h89 == io_inputs_1[7:0] ? 7'h0 : _GEN_5512; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5514 = 8'h8a == io_inputs_1[7:0] ? 7'h0 : _GEN_5513; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5515 = 8'h8b == io_inputs_1[7:0] ? 7'h0 : _GEN_5514; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5516 = 8'h8c == io_inputs_1[7:0] ? 7'h0 : _GEN_5515; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5517 = 8'h8d == io_inputs_1[7:0] ? 7'h0 : _GEN_5516; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5518 = 8'h8e == io_inputs_1[7:0] ? 7'h0 : _GEN_5517; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5519 = 8'h8f == io_inputs_1[7:0] ? 7'h0 : _GEN_5518; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5520 = 8'h90 == io_inputs_1[7:0] ? 7'h0 : _GEN_5519; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5521 = 8'h91 == io_inputs_1[7:0] ? 7'h0 : _GEN_5520; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5522 = 8'h92 == io_inputs_1[7:0] ? 7'h0 : _GEN_5521; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5523 = 8'h93 == io_inputs_1[7:0] ? 7'h0 : _GEN_5522; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5524 = 8'h94 == io_inputs_1[7:0] ? 7'h0 : _GEN_5523; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5525 = 8'h95 == io_inputs_1[7:0] ? 7'h0 : _GEN_5524; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5526 = 8'h96 == io_inputs_1[7:0] ? 7'h0 : _GEN_5525; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5527 = 8'h97 == io_inputs_1[7:0] ? 7'h0 : _GEN_5526; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5528 = 8'h98 == io_inputs_1[7:0] ? 7'h0 : _GEN_5527; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5529 = 8'h99 == io_inputs_1[7:0] ? 7'h0 : _GEN_5528; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5530 = 8'h9a == io_inputs_1[7:0] ? 7'h0 : _GEN_5529; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5531 = 8'h9b == io_inputs_1[7:0] ? 7'h0 : _GEN_5530; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5532 = 8'h9c == io_inputs_1[7:0] ? 7'h0 : _GEN_5531; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5533 = 8'h9d == io_inputs_1[7:0] ? 7'h0 : _GEN_5532; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5534 = 8'h9e == io_inputs_1[7:0] ? 7'h0 : _GEN_5533; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5535 = 8'h9f == io_inputs_1[7:0] ? 7'h0 : _GEN_5534; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5536 = 8'ha0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5535; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5537 = 8'ha1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5536; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5538 = 8'ha2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5537; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5539 = 8'ha3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5538; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5540 = 8'ha4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5539; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5541 = 8'ha5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5540; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5542 = 8'ha6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5541; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5543 = 8'ha7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5542; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5544 = 8'ha8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5543; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5545 = 8'ha9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5544; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5546 = 8'haa == io_inputs_1[7:0] ? 7'h0 : _GEN_5545; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5547 = 8'hab == io_inputs_1[7:0] ? 7'h0 : _GEN_5546; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5548 = 8'hac == io_inputs_1[7:0] ? 7'h0 : _GEN_5547; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5549 = 8'had == io_inputs_1[7:0] ? 7'h0 : _GEN_5548; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5550 = 8'hae == io_inputs_1[7:0] ? 7'h0 : _GEN_5549; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5551 = 8'haf == io_inputs_1[7:0] ? 7'h0 : _GEN_5550; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5552 = 8'hb0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5551; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5553 = 8'hb1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5552; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5554 = 8'hb2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5553; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5555 = 8'hb3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5554; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5556 = 8'hb4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5555; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5557 = 8'hb5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5556; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5558 = 8'hb6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5557; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5559 = 8'hb7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5558; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5560 = 8'hb8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5559; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5561 = 8'hb9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5560; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5562 = 8'hba == io_inputs_1[7:0] ? 7'h0 : _GEN_5561; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5563 = 8'hbb == io_inputs_1[7:0] ? 7'h0 : _GEN_5562; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5564 = 8'hbc == io_inputs_1[7:0] ? 7'h0 : _GEN_5563; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5565 = 8'hbd == io_inputs_1[7:0] ? 7'h0 : _GEN_5564; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5566 = 8'hbe == io_inputs_1[7:0] ? 7'h0 : _GEN_5565; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5567 = 8'hbf == io_inputs_1[7:0] ? 7'h0 : _GEN_5566; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5568 = 8'hc0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5567; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5569 = 8'hc1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5568; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5570 = 8'hc2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5569; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5571 = 8'hc3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5570; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5572 = 8'hc4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5571; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5573 = 8'hc5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5572; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5574 = 8'hc6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5573; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5575 = 8'hc7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5574; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5576 = 8'hc8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5575; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5577 = 8'hc9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5576; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5578 = 8'hca == io_inputs_1[7:0] ? 7'h0 : _GEN_5577; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5579 = 8'hcb == io_inputs_1[7:0] ? 7'h0 : _GEN_5578; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5580 = 8'hcc == io_inputs_1[7:0] ? 7'h0 : _GEN_5579; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5581 = 8'hcd == io_inputs_1[7:0] ? 7'h0 : _GEN_5580; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5582 = 8'hce == io_inputs_1[7:0] ? 7'h0 : _GEN_5581; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5583 = 8'hcf == io_inputs_1[7:0] ? 7'h0 : _GEN_5582; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5584 = 8'hd0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5583; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5585 = 8'hd1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5584; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5586 = 8'hd2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5585; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5587 = 8'hd3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5586; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5588 = 8'hd4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5587; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5589 = 8'hd5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5588; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5590 = 8'hd6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5589; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5591 = 8'hd7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5590; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5592 = 8'hd8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5591; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5593 = 8'hd9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5592; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5594 = 8'hda == io_inputs_1[7:0] ? 7'h0 : _GEN_5593; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5595 = 8'hdb == io_inputs_1[7:0] ? 7'h0 : _GEN_5594; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5596 = 8'hdc == io_inputs_1[7:0] ? 7'h0 : _GEN_5595; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5597 = 8'hdd == io_inputs_1[7:0] ? 7'h0 : _GEN_5596; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5598 = 8'hde == io_inputs_1[7:0] ? 7'h0 : _GEN_5597; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5599 = 8'hdf == io_inputs_1[7:0] ? 7'h0 : _GEN_5598; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5600 = 8'he0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5599; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5601 = 8'he1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5600; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5602 = 8'he2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5601; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5603 = 8'he3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5602; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5604 = 8'he4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5603; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5605 = 8'he5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5604; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5606 = 8'he6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5605; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5607 = 8'he7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5606; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5608 = 8'he8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5607; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5609 = 8'he9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5608; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5610 = 8'hea == io_inputs_1[7:0] ? 7'h0 : _GEN_5609; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5611 = 8'heb == io_inputs_1[7:0] ? 7'h0 : _GEN_5610; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5612 = 8'hec == io_inputs_1[7:0] ? 7'h0 : _GEN_5611; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5613 = 8'hed == io_inputs_1[7:0] ? 7'h0 : _GEN_5612; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5614 = 8'hee == io_inputs_1[7:0] ? 7'h0 : _GEN_5613; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5615 = 8'hef == io_inputs_1[7:0] ? 7'h0 : _GEN_5614; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5616 = 8'hf0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5615; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5617 = 8'hf1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5616; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5618 = 8'hf2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5617; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5619 = 8'hf3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5618; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5620 = 8'hf4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5619; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5621 = 8'hf5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5620; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5622 = 8'hf6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5621; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5623 = 8'hf7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5622; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5624 = 8'hf8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5623; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5625 = 8'hf9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5624; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5626 = 8'hfa == io_inputs_1[7:0] ? 7'h0 : _GEN_5625; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5627 = 8'hfb == io_inputs_1[7:0] ? 7'h0 : _GEN_5626; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5628 = 8'hfc == io_inputs_1[7:0] ? 7'h0 : _GEN_5627; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5693 = 8'h3d == io_inputs_1[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5694 = 8'h3e == io_inputs_1[7:0] ? 7'ha : _GEN_5693; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5695 = 8'h3f == io_inputs_1[7:0] ? 7'hf : _GEN_5694; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5696 = 8'h40 == io_inputs_1[7:0] ? 7'h14 : _GEN_5695; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5697 = 8'h41 == io_inputs_1[7:0] ? 7'h19 : _GEN_5696; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5698 = 8'h42 == io_inputs_1[7:0] ? 7'h1e : _GEN_5697; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5699 = 8'h43 == io_inputs_1[7:0] ? 7'h23 : _GEN_5698; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5700 = 8'h44 == io_inputs_1[7:0] ? 7'h28 : _GEN_5699; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5701 = 8'h45 == io_inputs_1[7:0] ? 7'h2d : _GEN_5700; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5702 = 8'h46 == io_inputs_1[7:0] ? 7'h32 : _GEN_5701; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5703 = 8'h47 == io_inputs_1[7:0] ? 7'h37 : _GEN_5702; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5704 = 8'h48 == io_inputs_1[7:0] ? 7'h3c : _GEN_5703; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5705 = 8'h49 == io_inputs_1[7:0] ? 7'h41 : _GEN_5704; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5706 = 8'h4a == io_inputs_1[7:0] ? 7'h46 : _GEN_5705; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5707 = 8'h4b == io_inputs_1[7:0] ? 7'h4b : _GEN_5706; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5708 = 8'h4c == io_inputs_1[7:0] ? 7'h50 : _GEN_5707; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5709 = 8'h4d == io_inputs_1[7:0] ? 7'h55 : _GEN_5708; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5710 = 8'h4e == io_inputs_1[7:0] ? 7'h5a : _GEN_5709; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5711 = 8'h4f == io_inputs_1[7:0] ? 7'h5f : _GEN_5710; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5712 = 8'h50 == io_inputs_1[7:0] ? 7'h64 : _GEN_5711; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5713 = 8'h51 == io_inputs_1[7:0] ? 7'h64 : _GEN_5712; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5714 = 8'h52 == io_inputs_1[7:0] ? 7'h64 : _GEN_5713; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5715 = 8'h53 == io_inputs_1[7:0] ? 7'h64 : _GEN_5714; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5716 = 8'h54 == io_inputs_1[7:0] ? 7'h64 : _GEN_5715; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5717 = 8'h55 == io_inputs_1[7:0] ? 7'h64 : _GEN_5716; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5718 = 8'h56 == io_inputs_1[7:0] ? 7'h64 : _GEN_5717; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5719 = 8'h57 == io_inputs_1[7:0] ? 7'h64 : _GEN_5718; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5720 = 8'h58 == io_inputs_1[7:0] ? 7'h64 : _GEN_5719; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5721 = 8'h59 == io_inputs_1[7:0] ? 7'h64 : _GEN_5720; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5722 = 8'h5a == io_inputs_1[7:0] ? 7'h64 : _GEN_5721; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5723 = 8'h5b == io_inputs_1[7:0] ? 7'h64 : _GEN_5722; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5724 = 8'h5c == io_inputs_1[7:0] ? 7'h64 : _GEN_5723; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5725 = 8'h5d == io_inputs_1[7:0] ? 7'h64 : _GEN_5724; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5726 = 8'h5e == io_inputs_1[7:0] ? 7'h64 : _GEN_5725; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5727 = 8'h5f == io_inputs_1[7:0] ? 7'h64 : _GEN_5726; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5728 = 8'h60 == io_inputs_1[7:0] ? 7'h64 : _GEN_5727; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5729 = 8'h61 == io_inputs_1[7:0] ? 7'h64 : _GEN_5728; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5730 = 8'h62 == io_inputs_1[7:0] ? 7'h64 : _GEN_5729; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5731 = 8'h63 == io_inputs_1[7:0] ? 7'h64 : _GEN_5730; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5732 = 8'h64 == io_inputs_1[7:0] ? 7'h64 : _GEN_5731; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5733 = 8'h65 == io_inputs_1[7:0] ? 7'h5f : _GEN_5732; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5734 = 8'h66 == io_inputs_1[7:0] ? 7'h5a : _GEN_5733; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5735 = 8'h67 == io_inputs_1[7:0] ? 7'h55 : _GEN_5734; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5736 = 8'h68 == io_inputs_1[7:0] ? 7'h50 : _GEN_5735; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5737 = 8'h69 == io_inputs_1[7:0] ? 7'h4b : _GEN_5736; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5738 = 8'h6a == io_inputs_1[7:0] ? 7'h46 : _GEN_5737; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5739 = 8'h6b == io_inputs_1[7:0] ? 7'h41 : _GEN_5738; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5740 = 8'h6c == io_inputs_1[7:0] ? 7'h3c : _GEN_5739; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5741 = 8'h6d == io_inputs_1[7:0] ? 7'h37 : _GEN_5740; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5742 = 8'h6e == io_inputs_1[7:0] ? 7'h32 : _GEN_5741; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5743 = 8'h6f == io_inputs_1[7:0] ? 7'h2d : _GEN_5742; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5744 = 8'h70 == io_inputs_1[7:0] ? 7'h28 : _GEN_5743; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5745 = 8'h71 == io_inputs_1[7:0] ? 7'h23 : _GEN_5744; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5746 = 8'h72 == io_inputs_1[7:0] ? 7'h1e : _GEN_5745; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5747 = 8'h73 == io_inputs_1[7:0] ? 7'h19 : _GEN_5746; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5748 = 8'h74 == io_inputs_1[7:0] ? 7'h14 : _GEN_5747; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5749 = 8'h75 == io_inputs_1[7:0] ? 7'hf : _GEN_5748; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5750 = 8'h76 == io_inputs_1[7:0] ? 7'ha : _GEN_5749; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5751 = 8'h77 == io_inputs_1[7:0] ? 7'h5 : _GEN_5750; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5752 = 8'h78 == io_inputs_1[7:0] ? 7'h0 : _GEN_5751; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5753 = 8'h79 == io_inputs_1[7:0] ? 7'h0 : _GEN_5752; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5754 = 8'h7a == io_inputs_1[7:0] ? 7'h0 : _GEN_5753; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5755 = 8'h7b == io_inputs_1[7:0] ? 7'h0 : _GEN_5754; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5756 = 8'h7c == io_inputs_1[7:0] ? 7'h0 : _GEN_5755; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5757 = 8'h7d == io_inputs_1[7:0] ? 7'h0 : _GEN_5756; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5758 = 8'h7e == io_inputs_1[7:0] ? 7'h0 : _GEN_5757; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5759 = 8'h7f == io_inputs_1[7:0] ? 7'h0 : _GEN_5758; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5760 = 8'h80 == io_inputs_1[7:0] ? 7'h0 : _GEN_5759; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5761 = 8'h81 == io_inputs_1[7:0] ? 7'h0 : _GEN_5760; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5762 = 8'h82 == io_inputs_1[7:0] ? 7'h0 : _GEN_5761; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5763 = 8'h83 == io_inputs_1[7:0] ? 7'h0 : _GEN_5762; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5764 = 8'h84 == io_inputs_1[7:0] ? 7'h0 : _GEN_5763; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5765 = 8'h85 == io_inputs_1[7:0] ? 7'h0 : _GEN_5764; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5766 = 8'h86 == io_inputs_1[7:0] ? 7'h0 : _GEN_5765; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5767 = 8'h87 == io_inputs_1[7:0] ? 7'h0 : _GEN_5766; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5768 = 8'h88 == io_inputs_1[7:0] ? 7'h0 : _GEN_5767; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5769 = 8'h89 == io_inputs_1[7:0] ? 7'h0 : _GEN_5768; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5770 = 8'h8a == io_inputs_1[7:0] ? 7'h0 : _GEN_5769; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5771 = 8'h8b == io_inputs_1[7:0] ? 7'h0 : _GEN_5770; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5772 = 8'h8c == io_inputs_1[7:0] ? 7'h0 : _GEN_5771; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5773 = 8'h8d == io_inputs_1[7:0] ? 7'h0 : _GEN_5772; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5774 = 8'h8e == io_inputs_1[7:0] ? 7'h0 : _GEN_5773; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5775 = 8'h8f == io_inputs_1[7:0] ? 7'h0 : _GEN_5774; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5776 = 8'h90 == io_inputs_1[7:0] ? 7'h0 : _GEN_5775; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5777 = 8'h91 == io_inputs_1[7:0] ? 7'h0 : _GEN_5776; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5778 = 8'h92 == io_inputs_1[7:0] ? 7'h0 : _GEN_5777; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5779 = 8'h93 == io_inputs_1[7:0] ? 7'h0 : _GEN_5778; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5780 = 8'h94 == io_inputs_1[7:0] ? 7'h0 : _GEN_5779; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5781 = 8'h95 == io_inputs_1[7:0] ? 7'h0 : _GEN_5780; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5782 = 8'h96 == io_inputs_1[7:0] ? 7'h0 : _GEN_5781; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5783 = 8'h97 == io_inputs_1[7:0] ? 7'h0 : _GEN_5782; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5784 = 8'h98 == io_inputs_1[7:0] ? 7'h0 : _GEN_5783; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5785 = 8'h99 == io_inputs_1[7:0] ? 7'h0 : _GEN_5784; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5786 = 8'h9a == io_inputs_1[7:0] ? 7'h0 : _GEN_5785; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5787 = 8'h9b == io_inputs_1[7:0] ? 7'h0 : _GEN_5786; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5788 = 8'h9c == io_inputs_1[7:0] ? 7'h0 : _GEN_5787; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5789 = 8'h9d == io_inputs_1[7:0] ? 7'h0 : _GEN_5788; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5790 = 8'h9e == io_inputs_1[7:0] ? 7'h0 : _GEN_5789; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5791 = 8'h9f == io_inputs_1[7:0] ? 7'h0 : _GEN_5790; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5792 = 8'ha0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5791; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5793 = 8'ha1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5792; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5794 = 8'ha2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5793; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5795 = 8'ha3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5794; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5796 = 8'ha4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5795; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5797 = 8'ha5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5796; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5798 = 8'ha6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5797; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5799 = 8'ha7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5798; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5800 = 8'ha8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5799; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5801 = 8'ha9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5800; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5802 = 8'haa == io_inputs_1[7:0] ? 7'h0 : _GEN_5801; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5803 = 8'hab == io_inputs_1[7:0] ? 7'h0 : _GEN_5802; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5804 = 8'hac == io_inputs_1[7:0] ? 7'h0 : _GEN_5803; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5805 = 8'had == io_inputs_1[7:0] ? 7'h0 : _GEN_5804; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5806 = 8'hae == io_inputs_1[7:0] ? 7'h0 : _GEN_5805; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5807 = 8'haf == io_inputs_1[7:0] ? 7'h0 : _GEN_5806; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5808 = 8'hb0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5807; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5809 = 8'hb1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5808; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5810 = 8'hb2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5809; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5811 = 8'hb3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5810; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5812 = 8'hb4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5811; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5813 = 8'hb5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5812; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5814 = 8'hb6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5813; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5815 = 8'hb7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5814; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5816 = 8'hb8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5815; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5817 = 8'hb9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5816; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5818 = 8'hba == io_inputs_1[7:0] ? 7'h0 : _GEN_5817; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5819 = 8'hbb == io_inputs_1[7:0] ? 7'h0 : _GEN_5818; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5820 = 8'hbc == io_inputs_1[7:0] ? 7'h0 : _GEN_5819; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5821 = 8'hbd == io_inputs_1[7:0] ? 7'h0 : _GEN_5820; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5822 = 8'hbe == io_inputs_1[7:0] ? 7'h0 : _GEN_5821; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5823 = 8'hbf == io_inputs_1[7:0] ? 7'h0 : _GEN_5822; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5824 = 8'hc0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5823; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5825 = 8'hc1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5824; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5826 = 8'hc2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5825; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5827 = 8'hc3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5826; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5828 = 8'hc4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5827; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5829 = 8'hc5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5828; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5830 = 8'hc6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5829; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5831 = 8'hc7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5830; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5832 = 8'hc8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5831; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5833 = 8'hc9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5832; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5834 = 8'hca == io_inputs_1[7:0] ? 7'h0 : _GEN_5833; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5835 = 8'hcb == io_inputs_1[7:0] ? 7'h0 : _GEN_5834; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5836 = 8'hcc == io_inputs_1[7:0] ? 7'h0 : _GEN_5835; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5837 = 8'hcd == io_inputs_1[7:0] ? 7'h0 : _GEN_5836; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5838 = 8'hce == io_inputs_1[7:0] ? 7'h0 : _GEN_5837; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5839 = 8'hcf == io_inputs_1[7:0] ? 7'h0 : _GEN_5838; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5840 = 8'hd0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5839; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5841 = 8'hd1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5840; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5842 = 8'hd2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5841; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5843 = 8'hd3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5842; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5844 = 8'hd4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5843; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5845 = 8'hd5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5844; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5846 = 8'hd6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5845; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5847 = 8'hd7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5846; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5848 = 8'hd8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5847; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5849 = 8'hd9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5848; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5850 = 8'hda == io_inputs_1[7:0] ? 7'h0 : _GEN_5849; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5851 = 8'hdb == io_inputs_1[7:0] ? 7'h0 : _GEN_5850; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5852 = 8'hdc == io_inputs_1[7:0] ? 7'h0 : _GEN_5851; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5853 = 8'hdd == io_inputs_1[7:0] ? 7'h0 : _GEN_5852; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5854 = 8'hde == io_inputs_1[7:0] ? 7'h0 : _GEN_5853; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5855 = 8'hdf == io_inputs_1[7:0] ? 7'h0 : _GEN_5854; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5856 = 8'he0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5855; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5857 = 8'he1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5856; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5858 = 8'he2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5857; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5859 = 8'he3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5858; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5860 = 8'he4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5859; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5861 = 8'he5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5860; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5862 = 8'he6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5861; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5863 = 8'he7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5862; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5864 = 8'he8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5863; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5865 = 8'he9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5864; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5866 = 8'hea == io_inputs_1[7:0] ? 7'h0 : _GEN_5865; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5867 = 8'heb == io_inputs_1[7:0] ? 7'h0 : _GEN_5866; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5868 = 8'hec == io_inputs_1[7:0] ? 7'h0 : _GEN_5867; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5869 = 8'hed == io_inputs_1[7:0] ? 7'h0 : _GEN_5868; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5870 = 8'hee == io_inputs_1[7:0] ? 7'h0 : _GEN_5869; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5871 = 8'hef == io_inputs_1[7:0] ? 7'h0 : _GEN_5870; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5872 = 8'hf0 == io_inputs_1[7:0] ? 7'h0 : _GEN_5871; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5873 = 8'hf1 == io_inputs_1[7:0] ? 7'h0 : _GEN_5872; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5874 = 8'hf2 == io_inputs_1[7:0] ? 7'h0 : _GEN_5873; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5875 = 8'hf3 == io_inputs_1[7:0] ? 7'h0 : _GEN_5874; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5876 = 8'hf4 == io_inputs_1[7:0] ? 7'h0 : _GEN_5875; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5877 = 8'hf5 == io_inputs_1[7:0] ? 7'h0 : _GEN_5876; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5878 = 8'hf6 == io_inputs_1[7:0] ? 7'h0 : _GEN_5877; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5879 = 8'hf7 == io_inputs_1[7:0] ? 7'h0 : _GEN_5878; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5880 = 8'hf8 == io_inputs_1[7:0] ? 7'h0 : _GEN_5879; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5881 = 8'hf9 == io_inputs_1[7:0] ? 7'h0 : _GEN_5880; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5882 = 8'hfa == io_inputs_1[7:0] ? 7'h0 : _GEN_5881; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5883 = 8'hfb == io_inputs_1[7:0] ? 7'h0 : _GEN_5882; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5884 = 8'hfc == io_inputs_1[7:0] ? 7'h0 : _GEN_5883; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5989 = 8'h65 == io_inputs_1[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5990 = 8'h66 == io_inputs_1[7:0] ? 7'ha : _GEN_5989; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5991 = 8'h67 == io_inputs_1[7:0] ? 7'hf : _GEN_5990; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5992 = 8'h68 == io_inputs_1[7:0] ? 7'h14 : _GEN_5991; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5993 = 8'h69 == io_inputs_1[7:0] ? 7'h19 : _GEN_5992; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5994 = 8'h6a == io_inputs_1[7:0] ? 7'h1e : _GEN_5993; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5995 = 8'h6b == io_inputs_1[7:0] ? 7'h23 : _GEN_5994; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5996 = 8'h6c == io_inputs_1[7:0] ? 7'h28 : _GEN_5995; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5997 = 8'h6d == io_inputs_1[7:0] ? 7'h2d : _GEN_5996; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5998 = 8'h6e == io_inputs_1[7:0] ? 7'h32 : _GEN_5997; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_5999 = 8'h6f == io_inputs_1[7:0] ? 7'h37 : _GEN_5998; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6000 = 8'h70 == io_inputs_1[7:0] ? 7'h3c : _GEN_5999; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6001 = 8'h71 == io_inputs_1[7:0] ? 7'h41 : _GEN_6000; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6002 = 8'h72 == io_inputs_1[7:0] ? 7'h46 : _GEN_6001; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6003 = 8'h73 == io_inputs_1[7:0] ? 7'h4b : _GEN_6002; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6004 = 8'h74 == io_inputs_1[7:0] ? 7'h50 : _GEN_6003; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6005 = 8'h75 == io_inputs_1[7:0] ? 7'h55 : _GEN_6004; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6006 = 8'h76 == io_inputs_1[7:0] ? 7'h5a : _GEN_6005; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6007 = 8'h77 == io_inputs_1[7:0] ? 7'h5f : _GEN_6006; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6008 = 8'h78 == io_inputs_1[7:0] ? 7'h64 : _GEN_6007; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6009 = 8'h79 == io_inputs_1[7:0] ? 7'h64 : _GEN_6008; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6010 = 8'h7a == io_inputs_1[7:0] ? 7'h64 : _GEN_6009; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6011 = 8'h7b == io_inputs_1[7:0] ? 7'h64 : _GEN_6010; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6012 = 8'h7c == io_inputs_1[7:0] ? 7'h64 : _GEN_6011; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6013 = 8'h7d == io_inputs_1[7:0] ? 7'h64 : _GEN_6012; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6014 = 8'h7e == io_inputs_1[7:0] ? 7'h64 : _GEN_6013; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6015 = 8'h7f == io_inputs_1[7:0] ? 7'h64 : _GEN_6014; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6016 = 8'h80 == io_inputs_1[7:0] ? 7'h64 : _GEN_6015; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6017 = 8'h81 == io_inputs_1[7:0] ? 7'h64 : _GEN_6016; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6018 = 8'h82 == io_inputs_1[7:0] ? 7'h64 : _GEN_6017; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6019 = 8'h83 == io_inputs_1[7:0] ? 7'h64 : _GEN_6018; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6020 = 8'h84 == io_inputs_1[7:0] ? 7'h64 : _GEN_6019; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6021 = 8'h85 == io_inputs_1[7:0] ? 7'h64 : _GEN_6020; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6022 = 8'h86 == io_inputs_1[7:0] ? 7'h64 : _GEN_6021; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6023 = 8'h87 == io_inputs_1[7:0] ? 7'h64 : _GEN_6022; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6024 = 8'h88 == io_inputs_1[7:0] ? 7'h64 : _GEN_6023; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6025 = 8'h89 == io_inputs_1[7:0] ? 7'h64 : _GEN_6024; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6026 = 8'h8a == io_inputs_1[7:0] ? 7'h64 : _GEN_6025; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6027 = 8'h8b == io_inputs_1[7:0] ? 7'h64 : _GEN_6026; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6028 = 8'h8c == io_inputs_1[7:0] ? 7'h64 : _GEN_6027; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6029 = 8'h8d == io_inputs_1[7:0] ? 7'h5f : _GEN_6028; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6030 = 8'h8e == io_inputs_1[7:0] ? 7'h5a : _GEN_6029; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6031 = 8'h8f == io_inputs_1[7:0] ? 7'h55 : _GEN_6030; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6032 = 8'h90 == io_inputs_1[7:0] ? 7'h50 : _GEN_6031; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6033 = 8'h91 == io_inputs_1[7:0] ? 7'h4b : _GEN_6032; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6034 = 8'h92 == io_inputs_1[7:0] ? 7'h46 : _GEN_6033; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6035 = 8'h93 == io_inputs_1[7:0] ? 7'h41 : _GEN_6034; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6036 = 8'h94 == io_inputs_1[7:0] ? 7'h3c : _GEN_6035; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6037 = 8'h95 == io_inputs_1[7:0] ? 7'h37 : _GEN_6036; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6038 = 8'h96 == io_inputs_1[7:0] ? 7'h32 : _GEN_6037; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6039 = 8'h97 == io_inputs_1[7:0] ? 7'h2d : _GEN_6038; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6040 = 8'h98 == io_inputs_1[7:0] ? 7'h28 : _GEN_6039; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6041 = 8'h99 == io_inputs_1[7:0] ? 7'h23 : _GEN_6040; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6042 = 8'h9a == io_inputs_1[7:0] ? 7'h1e : _GEN_6041; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6043 = 8'h9b == io_inputs_1[7:0] ? 7'h19 : _GEN_6042; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6044 = 8'h9c == io_inputs_1[7:0] ? 7'h14 : _GEN_6043; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6045 = 8'h9d == io_inputs_1[7:0] ? 7'hf : _GEN_6044; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6046 = 8'h9e == io_inputs_1[7:0] ? 7'ha : _GEN_6045; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6047 = 8'h9f == io_inputs_1[7:0] ? 7'h5 : _GEN_6046; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6048 = 8'ha0 == io_inputs_1[7:0] ? 7'h0 : _GEN_6047; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6049 = 8'ha1 == io_inputs_1[7:0] ? 7'h0 : _GEN_6048; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6050 = 8'ha2 == io_inputs_1[7:0] ? 7'h0 : _GEN_6049; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6051 = 8'ha3 == io_inputs_1[7:0] ? 7'h0 : _GEN_6050; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6052 = 8'ha4 == io_inputs_1[7:0] ? 7'h0 : _GEN_6051; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6053 = 8'ha5 == io_inputs_1[7:0] ? 7'h0 : _GEN_6052; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6054 = 8'ha6 == io_inputs_1[7:0] ? 7'h0 : _GEN_6053; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6055 = 8'ha7 == io_inputs_1[7:0] ? 7'h0 : _GEN_6054; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6056 = 8'ha8 == io_inputs_1[7:0] ? 7'h0 : _GEN_6055; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6057 = 8'ha9 == io_inputs_1[7:0] ? 7'h0 : _GEN_6056; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6058 = 8'haa == io_inputs_1[7:0] ? 7'h0 : _GEN_6057; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6059 = 8'hab == io_inputs_1[7:0] ? 7'h0 : _GEN_6058; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6060 = 8'hac == io_inputs_1[7:0] ? 7'h0 : _GEN_6059; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6061 = 8'had == io_inputs_1[7:0] ? 7'h0 : _GEN_6060; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6062 = 8'hae == io_inputs_1[7:0] ? 7'h0 : _GEN_6061; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6063 = 8'haf == io_inputs_1[7:0] ? 7'h0 : _GEN_6062; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6064 = 8'hb0 == io_inputs_1[7:0] ? 7'h0 : _GEN_6063; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6065 = 8'hb1 == io_inputs_1[7:0] ? 7'h0 : _GEN_6064; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6066 = 8'hb2 == io_inputs_1[7:0] ? 7'h0 : _GEN_6065; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6067 = 8'hb3 == io_inputs_1[7:0] ? 7'h0 : _GEN_6066; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6068 = 8'hb4 == io_inputs_1[7:0] ? 7'h0 : _GEN_6067; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6069 = 8'hb5 == io_inputs_1[7:0] ? 7'h0 : _GEN_6068; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6070 = 8'hb6 == io_inputs_1[7:0] ? 7'h0 : _GEN_6069; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6071 = 8'hb7 == io_inputs_1[7:0] ? 7'h0 : _GEN_6070; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6072 = 8'hb8 == io_inputs_1[7:0] ? 7'h0 : _GEN_6071; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6073 = 8'hb9 == io_inputs_1[7:0] ? 7'h0 : _GEN_6072; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6074 = 8'hba == io_inputs_1[7:0] ? 7'h0 : _GEN_6073; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6075 = 8'hbb == io_inputs_1[7:0] ? 7'h0 : _GEN_6074; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6076 = 8'hbc == io_inputs_1[7:0] ? 7'h0 : _GEN_6075; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6077 = 8'hbd == io_inputs_1[7:0] ? 7'h0 : _GEN_6076; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6078 = 8'hbe == io_inputs_1[7:0] ? 7'h0 : _GEN_6077; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6079 = 8'hbf == io_inputs_1[7:0] ? 7'h0 : _GEN_6078; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6080 = 8'hc0 == io_inputs_1[7:0] ? 7'h0 : _GEN_6079; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6081 = 8'hc1 == io_inputs_1[7:0] ? 7'h0 : _GEN_6080; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6082 = 8'hc2 == io_inputs_1[7:0] ? 7'h0 : _GEN_6081; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6083 = 8'hc3 == io_inputs_1[7:0] ? 7'h0 : _GEN_6082; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6084 = 8'hc4 == io_inputs_1[7:0] ? 7'h0 : _GEN_6083; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6085 = 8'hc5 == io_inputs_1[7:0] ? 7'h0 : _GEN_6084; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6086 = 8'hc6 == io_inputs_1[7:0] ? 7'h0 : _GEN_6085; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6087 = 8'hc7 == io_inputs_1[7:0] ? 7'h0 : _GEN_6086; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6088 = 8'hc8 == io_inputs_1[7:0] ? 7'h0 : _GEN_6087; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6089 = 8'hc9 == io_inputs_1[7:0] ? 7'h0 : _GEN_6088; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6090 = 8'hca == io_inputs_1[7:0] ? 7'h0 : _GEN_6089; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6091 = 8'hcb == io_inputs_1[7:0] ? 7'h0 : _GEN_6090; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6092 = 8'hcc == io_inputs_1[7:0] ? 7'h0 : _GEN_6091; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6093 = 8'hcd == io_inputs_1[7:0] ? 7'h0 : _GEN_6092; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6094 = 8'hce == io_inputs_1[7:0] ? 7'h0 : _GEN_6093; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6095 = 8'hcf == io_inputs_1[7:0] ? 7'h0 : _GEN_6094; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6096 = 8'hd0 == io_inputs_1[7:0] ? 7'h0 : _GEN_6095; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6097 = 8'hd1 == io_inputs_1[7:0] ? 7'h0 : _GEN_6096; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6098 = 8'hd2 == io_inputs_1[7:0] ? 7'h0 : _GEN_6097; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6099 = 8'hd3 == io_inputs_1[7:0] ? 7'h0 : _GEN_6098; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6100 = 8'hd4 == io_inputs_1[7:0] ? 7'h0 : _GEN_6099; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6101 = 8'hd5 == io_inputs_1[7:0] ? 7'h0 : _GEN_6100; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6102 = 8'hd6 == io_inputs_1[7:0] ? 7'h0 : _GEN_6101; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6103 = 8'hd7 == io_inputs_1[7:0] ? 7'h0 : _GEN_6102; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6104 = 8'hd8 == io_inputs_1[7:0] ? 7'h0 : _GEN_6103; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6105 = 8'hd9 == io_inputs_1[7:0] ? 7'h0 : _GEN_6104; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6106 = 8'hda == io_inputs_1[7:0] ? 7'h0 : _GEN_6105; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6107 = 8'hdb == io_inputs_1[7:0] ? 7'h0 : _GEN_6106; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6108 = 8'hdc == io_inputs_1[7:0] ? 7'h0 : _GEN_6107; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6109 = 8'hdd == io_inputs_1[7:0] ? 7'h0 : _GEN_6108; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6110 = 8'hde == io_inputs_1[7:0] ? 7'h0 : _GEN_6109; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6111 = 8'hdf == io_inputs_1[7:0] ? 7'h0 : _GEN_6110; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6112 = 8'he0 == io_inputs_1[7:0] ? 7'h0 : _GEN_6111; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6113 = 8'he1 == io_inputs_1[7:0] ? 7'h0 : _GEN_6112; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6114 = 8'he2 == io_inputs_1[7:0] ? 7'h0 : _GEN_6113; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6115 = 8'he3 == io_inputs_1[7:0] ? 7'h0 : _GEN_6114; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6116 = 8'he4 == io_inputs_1[7:0] ? 7'h0 : _GEN_6115; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6117 = 8'he5 == io_inputs_1[7:0] ? 7'h0 : _GEN_6116; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6118 = 8'he6 == io_inputs_1[7:0] ? 7'h0 : _GEN_6117; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6119 = 8'he7 == io_inputs_1[7:0] ? 7'h0 : _GEN_6118; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6120 = 8'he8 == io_inputs_1[7:0] ? 7'h0 : _GEN_6119; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6121 = 8'he9 == io_inputs_1[7:0] ? 7'h0 : _GEN_6120; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6122 = 8'hea == io_inputs_1[7:0] ? 7'h0 : _GEN_6121; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6123 = 8'heb == io_inputs_1[7:0] ? 7'h0 : _GEN_6122; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6124 = 8'hec == io_inputs_1[7:0] ? 7'h0 : _GEN_6123; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6125 = 8'hed == io_inputs_1[7:0] ? 7'h0 : _GEN_6124; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6126 = 8'hee == io_inputs_1[7:0] ? 7'h0 : _GEN_6125; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6127 = 8'hef == io_inputs_1[7:0] ? 7'h0 : _GEN_6126; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6128 = 8'hf0 == io_inputs_1[7:0] ? 7'h0 : _GEN_6127; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6129 = 8'hf1 == io_inputs_1[7:0] ? 7'h0 : _GEN_6128; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6130 = 8'hf2 == io_inputs_1[7:0] ? 7'h0 : _GEN_6129; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6131 = 8'hf3 == io_inputs_1[7:0] ? 7'h0 : _GEN_6130; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6132 = 8'hf4 == io_inputs_1[7:0] ? 7'h0 : _GEN_6131; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6133 = 8'hf5 == io_inputs_1[7:0] ? 7'h0 : _GEN_6132; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6134 = 8'hf6 == io_inputs_1[7:0] ? 7'h0 : _GEN_6133; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6135 = 8'hf7 == io_inputs_1[7:0] ? 7'h0 : _GEN_6134; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6136 = 8'hf8 == io_inputs_1[7:0] ? 7'h0 : _GEN_6135; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6137 = 8'hf9 == io_inputs_1[7:0] ? 7'h0 : _GEN_6136; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6138 = 8'hfa == io_inputs_1[7:0] ? 7'h0 : _GEN_6137; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6139 = 8'hfb == io_inputs_1[7:0] ? 7'h0 : _GEN_6138; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6140 = 8'hfc == io_inputs_1[7:0] ? 7'h0 : _GEN_6139; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6285 = 8'h8d == io_inputs_1[7:0] ? 7'h5 : 7'h0; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6286 = 8'h8e == io_inputs_1[7:0] ? 7'ha : _GEN_6285; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6287 = 8'h8f == io_inputs_1[7:0] ? 7'hf : _GEN_6286; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6288 = 8'h90 == io_inputs_1[7:0] ? 7'h14 : _GEN_6287; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6289 = 8'h91 == io_inputs_1[7:0] ? 7'h19 : _GEN_6288; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6290 = 8'h92 == io_inputs_1[7:0] ? 7'h1e : _GEN_6289; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6291 = 8'h93 == io_inputs_1[7:0] ? 7'h23 : _GEN_6290; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6292 = 8'h94 == io_inputs_1[7:0] ? 7'h28 : _GEN_6291; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6293 = 8'h95 == io_inputs_1[7:0] ? 7'h2d : _GEN_6292; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6294 = 8'h96 == io_inputs_1[7:0] ? 7'h32 : _GEN_6293; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6295 = 8'h97 == io_inputs_1[7:0] ? 7'h37 : _GEN_6294; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6296 = 8'h98 == io_inputs_1[7:0] ? 7'h3c : _GEN_6295; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6297 = 8'h99 == io_inputs_1[7:0] ? 7'h41 : _GEN_6296; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6298 = 8'h9a == io_inputs_1[7:0] ? 7'h46 : _GEN_6297; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6299 = 8'h9b == io_inputs_1[7:0] ? 7'h4b : _GEN_6298; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6300 = 8'h9c == io_inputs_1[7:0] ? 7'h50 : _GEN_6299; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6301 = 8'h9d == io_inputs_1[7:0] ? 7'h55 : _GEN_6300; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6302 = 8'h9e == io_inputs_1[7:0] ? 7'h5a : _GEN_6301; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6303 = 8'h9f == io_inputs_1[7:0] ? 7'h5f : _GEN_6302; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6304 = 8'ha0 == io_inputs_1[7:0] ? 7'h64 : _GEN_6303; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6305 = 8'ha1 == io_inputs_1[7:0] ? 7'h64 : _GEN_6304; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6306 = 8'ha2 == io_inputs_1[7:0] ? 7'h64 : _GEN_6305; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6307 = 8'ha3 == io_inputs_1[7:0] ? 7'h64 : _GEN_6306; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6308 = 8'ha4 == io_inputs_1[7:0] ? 7'h64 : _GEN_6307; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6309 = 8'ha5 == io_inputs_1[7:0] ? 7'h64 : _GEN_6308; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6310 = 8'ha6 == io_inputs_1[7:0] ? 7'h64 : _GEN_6309; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6311 = 8'ha7 == io_inputs_1[7:0] ? 7'h64 : _GEN_6310; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6312 = 8'ha8 == io_inputs_1[7:0] ? 7'h64 : _GEN_6311; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6313 = 8'ha9 == io_inputs_1[7:0] ? 7'h64 : _GEN_6312; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6314 = 8'haa == io_inputs_1[7:0] ? 7'h64 : _GEN_6313; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6315 = 8'hab == io_inputs_1[7:0] ? 7'h64 : _GEN_6314; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6316 = 8'hac == io_inputs_1[7:0] ? 7'h64 : _GEN_6315; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6317 = 8'had == io_inputs_1[7:0] ? 7'h64 : _GEN_6316; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6318 = 8'hae == io_inputs_1[7:0] ? 7'h64 : _GEN_6317; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6319 = 8'haf == io_inputs_1[7:0] ? 7'h64 : _GEN_6318; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6320 = 8'hb0 == io_inputs_1[7:0] ? 7'h64 : _GEN_6319; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6321 = 8'hb1 == io_inputs_1[7:0] ? 7'h64 : _GEN_6320; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6322 = 8'hb2 == io_inputs_1[7:0] ? 7'h64 : _GEN_6321; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6323 = 8'hb3 == io_inputs_1[7:0] ? 7'h64 : _GEN_6322; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6324 = 8'hb4 == io_inputs_1[7:0] ? 7'h64 : _GEN_6323; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6325 = 8'hb5 == io_inputs_1[7:0] ? 7'h64 : _GEN_6324; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6326 = 8'hb6 == io_inputs_1[7:0] ? 7'h64 : _GEN_6325; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6327 = 8'hb7 == io_inputs_1[7:0] ? 7'h64 : _GEN_6326; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6328 = 8'hb8 == io_inputs_1[7:0] ? 7'h64 : _GEN_6327; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6329 = 8'hb9 == io_inputs_1[7:0] ? 7'h64 : _GEN_6328; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6330 = 8'hba == io_inputs_1[7:0] ? 7'h64 : _GEN_6329; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6331 = 8'hbb == io_inputs_1[7:0] ? 7'h64 : _GEN_6330; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6332 = 8'hbc == io_inputs_1[7:0] ? 7'h64 : _GEN_6331; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6333 = 8'hbd == io_inputs_1[7:0] ? 7'h64 : _GEN_6332; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6334 = 8'hbe == io_inputs_1[7:0] ? 7'h64 : _GEN_6333; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6335 = 8'hbf == io_inputs_1[7:0] ? 7'h64 : _GEN_6334; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6336 = 8'hc0 == io_inputs_1[7:0] ? 7'h64 : _GEN_6335; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6337 = 8'hc1 == io_inputs_1[7:0] ? 7'h64 : _GEN_6336; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6338 = 8'hc2 == io_inputs_1[7:0] ? 7'h64 : _GEN_6337; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6339 = 8'hc3 == io_inputs_1[7:0] ? 7'h64 : _GEN_6338; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6340 = 8'hc4 == io_inputs_1[7:0] ? 7'h64 : _GEN_6339; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6341 = 8'hc5 == io_inputs_1[7:0] ? 7'h64 : _GEN_6340; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6342 = 8'hc6 == io_inputs_1[7:0] ? 7'h64 : _GEN_6341; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6343 = 8'hc7 == io_inputs_1[7:0] ? 7'h64 : _GEN_6342; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6344 = 8'hc8 == io_inputs_1[7:0] ? 7'h64 : _GEN_6343; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6345 = 8'hc9 == io_inputs_1[7:0] ? 7'h64 : _GEN_6344; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6346 = 8'hca == io_inputs_1[7:0] ? 7'h64 : _GEN_6345; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6347 = 8'hcb == io_inputs_1[7:0] ? 7'h64 : _GEN_6346; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6348 = 8'hcc == io_inputs_1[7:0] ? 7'h64 : _GEN_6347; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6349 = 8'hcd == io_inputs_1[7:0] ? 7'h64 : _GEN_6348; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6350 = 8'hce == io_inputs_1[7:0] ? 7'h64 : _GEN_6349; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6351 = 8'hcf == io_inputs_1[7:0] ? 7'h64 : _GEN_6350; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6352 = 8'hd0 == io_inputs_1[7:0] ? 7'h64 : _GEN_6351; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6353 = 8'hd1 == io_inputs_1[7:0] ? 7'h64 : _GEN_6352; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6354 = 8'hd2 == io_inputs_1[7:0] ? 7'h64 : _GEN_6353; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6355 = 8'hd3 == io_inputs_1[7:0] ? 7'h64 : _GEN_6354; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6356 = 8'hd4 == io_inputs_1[7:0] ? 7'h64 : _GEN_6355; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6357 = 8'hd5 == io_inputs_1[7:0] ? 7'h64 : _GEN_6356; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6358 = 8'hd6 == io_inputs_1[7:0] ? 7'h64 : _GEN_6357; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6359 = 8'hd7 == io_inputs_1[7:0] ? 7'h64 : _GEN_6358; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6360 = 8'hd8 == io_inputs_1[7:0] ? 7'h64 : _GEN_6359; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6361 = 8'hd9 == io_inputs_1[7:0] ? 7'h64 : _GEN_6360; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6362 = 8'hda == io_inputs_1[7:0] ? 7'h64 : _GEN_6361; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6363 = 8'hdb == io_inputs_1[7:0] ? 7'h64 : _GEN_6362; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6364 = 8'hdc == io_inputs_1[7:0] ? 7'h64 : _GEN_6363; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6365 = 8'hdd == io_inputs_1[7:0] ? 7'h64 : _GEN_6364; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6366 = 8'hde == io_inputs_1[7:0] ? 7'h64 : _GEN_6365; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6367 = 8'hdf == io_inputs_1[7:0] ? 7'h64 : _GEN_6366; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6368 = 8'he0 == io_inputs_1[7:0] ? 7'h64 : _GEN_6367; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6369 = 8'he1 == io_inputs_1[7:0] ? 7'h64 : _GEN_6368; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6370 = 8'he2 == io_inputs_1[7:0] ? 7'h64 : _GEN_6369; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6371 = 8'he3 == io_inputs_1[7:0] ? 7'h64 : _GEN_6370; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6372 = 8'he4 == io_inputs_1[7:0] ? 7'h64 : _GEN_6371; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6373 = 8'he5 == io_inputs_1[7:0] ? 7'h64 : _GEN_6372; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6374 = 8'he6 == io_inputs_1[7:0] ? 7'h64 : _GEN_6373; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6375 = 8'he7 == io_inputs_1[7:0] ? 7'h64 : _GEN_6374; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6376 = 8'he8 == io_inputs_1[7:0] ? 7'h64 : _GEN_6375; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6377 = 8'he9 == io_inputs_1[7:0] ? 7'h64 : _GEN_6376; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6378 = 8'hea == io_inputs_1[7:0] ? 7'h64 : _GEN_6377; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6379 = 8'heb == io_inputs_1[7:0] ? 7'h64 : _GEN_6378; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6380 = 8'hec == io_inputs_1[7:0] ? 7'h64 : _GEN_6379; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6381 = 8'hed == io_inputs_1[7:0] ? 7'h64 : _GEN_6380; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6382 = 8'hee == io_inputs_1[7:0] ? 7'h64 : _GEN_6381; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6383 = 8'hef == io_inputs_1[7:0] ? 7'h64 : _GEN_6382; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6384 = 8'hf0 == io_inputs_1[7:0] ? 7'h64 : _GEN_6383; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6385 = 8'hf1 == io_inputs_1[7:0] ? 7'h64 : _GEN_6384; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6386 = 8'hf2 == io_inputs_1[7:0] ? 7'h64 : _GEN_6385; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6387 = 8'hf3 == io_inputs_1[7:0] ? 7'h64 : _GEN_6386; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6388 = 8'hf4 == io_inputs_1[7:0] ? 7'h64 : _GEN_6387; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6389 = 8'hf5 == io_inputs_1[7:0] ? 7'h64 : _GEN_6388; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6390 = 8'hf6 == io_inputs_1[7:0] ? 7'h64 : _GEN_6389; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6391 = 8'hf7 == io_inputs_1[7:0] ? 7'h64 : _GEN_6390; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6392 = 8'hf8 == io_inputs_1[7:0] ? 7'h64 : _GEN_6391; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6393 = 8'hf9 == io_inputs_1[7:0] ? 7'h64 : _GEN_6392; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6394 = 8'hfa == io_inputs_1[7:0] ? 7'h64 : _GEN_6393; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6395 = 8'hfb == io_inputs_1[7:0] ? 7'h64 : _GEN_6394; // @[regular_fuzzification.scala 194:{38,38}]
  wire [6:0] _GEN_6396 = 8'hfc == io_inputs_1[7:0] ? 7'h64 : _GEN_6395; // @[regular_fuzzification.scala 194:{38,38}]
  wire  regMinVec_0_maxMinOutput = regMinVec_0_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_1_maxMinOutput = regMinVec_1_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_2_maxMinOutput = regMinVec_2_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_3_maxMinOutput = regMinVec_3_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_4_maxMinOutput = regMinVec_4_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_5_maxMinOutput = regMinVec_5_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_6_maxMinOutput = regMinVec_6_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_7_maxMinOutput = regMinVec_7_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_8_maxMinOutput = regMinVec_8_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_9_maxMinOutput = regMinVec_9_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_10_maxMinOutput = regMinVec_10_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_11_maxMinOutput = regMinVec_11_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_12_maxMinOutput = regMinVec_12_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_13_maxMinOutput = regMinVec_13_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_14_maxMinOutput = regMinVec_14_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_15_maxMinOutput = regMinVec_15_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_16_maxMinOutput = regMinVec_16_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_17_maxMinOutput = regMinVec_17_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_18_maxMinOutput = regMinVec_18_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_19_maxMinOutput = regMinVec_19_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_20_maxMinOutput = regMinVec_20_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_21_maxMinOutput = regMinVec_21_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_22_maxMinOutput = regMinVec_22_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_23_maxMinOutput = regMinVec_23_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire  regMinVec_24_maxMinOutput = regMinVec_24_comparatorModule_io_maxMin; // @[comparator.scala 71:28 90:18]
  wire [6:0] regMaxVec_0_result = regMaxVec_0_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [6:0] regMaxVec_1_result = regMaxVec_1_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [6:0] regMaxVec_2_result = regMaxVec_2_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [6:0] regMaxVec_3_result = regMaxVec_3_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [6:0] regMaxVec_4_result = regMaxVec_4_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  wire [6:0] outResult_result = outResult_comparatorModule_io_result; // @[multiple_comparator.scala 304:22 312:12]
  Comparator regMinVec_0_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_0_comparatorModule_io_in1),
    .io_in2(regMinVec_0_comparatorModule_io_in2),
    .io_maxMin(regMinVec_0_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_1_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_1_comparatorModule_io_in1),
    .io_in2(regMinVec_1_comparatorModule_io_in2),
    .io_maxMin(regMinVec_1_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_2_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_2_comparatorModule_io_in1),
    .io_in2(regMinVec_2_comparatorModule_io_in2),
    .io_maxMin(regMinVec_2_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_3_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_3_comparatorModule_io_in1),
    .io_in2(regMinVec_3_comparatorModule_io_in2),
    .io_maxMin(regMinVec_3_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_4_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_4_comparatorModule_io_in1),
    .io_in2(regMinVec_4_comparatorModule_io_in2),
    .io_maxMin(regMinVec_4_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_5_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_5_comparatorModule_io_in1),
    .io_in2(regMinVec_5_comparatorModule_io_in2),
    .io_maxMin(regMinVec_5_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_6_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_6_comparatorModule_io_in1),
    .io_in2(regMinVec_6_comparatorModule_io_in2),
    .io_maxMin(regMinVec_6_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_7_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_7_comparatorModule_io_in1),
    .io_in2(regMinVec_7_comparatorModule_io_in2),
    .io_maxMin(regMinVec_7_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_8_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_8_comparatorModule_io_in1),
    .io_in2(regMinVec_8_comparatorModule_io_in2),
    .io_maxMin(regMinVec_8_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_9_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_9_comparatorModule_io_in1),
    .io_in2(regMinVec_9_comparatorModule_io_in2),
    .io_maxMin(regMinVec_9_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_10_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_10_comparatorModule_io_in1),
    .io_in2(regMinVec_10_comparatorModule_io_in2),
    .io_maxMin(regMinVec_10_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_11_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_11_comparatorModule_io_in1),
    .io_in2(regMinVec_11_comparatorModule_io_in2),
    .io_maxMin(regMinVec_11_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_12_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_12_comparatorModule_io_in1),
    .io_in2(regMinVec_12_comparatorModule_io_in2),
    .io_maxMin(regMinVec_12_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_13_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_13_comparatorModule_io_in1),
    .io_in2(regMinVec_13_comparatorModule_io_in2),
    .io_maxMin(regMinVec_13_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_14_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_14_comparatorModule_io_in1),
    .io_in2(regMinVec_14_comparatorModule_io_in2),
    .io_maxMin(regMinVec_14_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_15_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_15_comparatorModule_io_in1),
    .io_in2(regMinVec_15_comparatorModule_io_in2),
    .io_maxMin(regMinVec_15_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_16_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_16_comparatorModule_io_in1),
    .io_in2(regMinVec_16_comparatorModule_io_in2),
    .io_maxMin(regMinVec_16_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_17_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_17_comparatorModule_io_in1),
    .io_in2(regMinVec_17_comparatorModule_io_in2),
    .io_maxMin(regMinVec_17_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_18_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_18_comparatorModule_io_in1),
    .io_in2(regMinVec_18_comparatorModule_io_in2),
    .io_maxMin(regMinVec_18_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_19_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_19_comparatorModule_io_in1),
    .io_in2(regMinVec_19_comparatorModule_io_in2),
    .io_maxMin(regMinVec_19_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_20_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_20_comparatorModule_io_in1),
    .io_in2(regMinVec_20_comparatorModule_io_in2),
    .io_maxMin(regMinVec_20_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_21_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_21_comparatorModule_io_in1),
    .io_in2(regMinVec_21_comparatorModule_io_in2),
    .io_maxMin(regMinVec_21_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_22_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_22_comparatorModule_io_in1),
    .io_in2(regMinVec_22_comparatorModule_io_in2),
    .io_maxMin(regMinVec_22_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_23_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_23_comparatorModule_io_in1),
    .io_in2(regMinVec_23_comparatorModule_io_in2),
    .io_maxMin(regMinVec_23_comparatorModule_io_maxMin)
  );
  Comparator regMinVec_24_comparatorModule ( // @[comparator.scala 69:34]
    .io_in1(regMinVec_24_comparatorModule_io_in1),
    .io_in2(regMinVec_24_comparatorModule_io_in2),
    .io_maxMin(regMinVec_24_comparatorModule_io_maxMin)
  );
  MultipleComparator regMaxVec_0_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_0_comparatorModule_clock),
    .io_start(regMaxVec_0_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_0_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_0_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_0_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_0_comparatorModule_io_inputs_3),
    .io_result(regMaxVec_0_comparatorModule_io_result)
  );
  MultipleComparator_1 regMaxVec_1_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_1_comparatorModule_clock),
    .io_start(regMaxVec_1_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_1_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_1_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_1_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_1_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_1_comparatorModule_io_inputs_4),
    .io_inputs_5(regMaxVec_1_comparatorModule_io_inputs_5),
    .io_result(regMaxVec_1_comparatorModule_io_result)
  );
  MultipleComparator regMaxVec_2_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_2_comparatorModule_clock),
    .io_start(regMaxVec_2_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_2_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_2_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_2_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_2_comparatorModule_io_inputs_3),
    .io_result(regMaxVec_2_comparatorModule_io_result)
  );
  MultipleComparator_1 regMaxVec_3_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_3_comparatorModule_clock),
    .io_start(regMaxVec_3_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_3_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_3_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_3_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_3_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_3_comparatorModule_io_inputs_4),
    .io_inputs_5(regMaxVec_3_comparatorModule_io_inputs_5),
    .io_result(regMaxVec_3_comparatorModule_io_result)
  );
  MultipleComparator_4 regMaxVec_4_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(regMaxVec_4_comparatorModule_clock),
    .io_start(regMaxVec_4_comparatorModule_io_start),
    .io_inputs_0(regMaxVec_4_comparatorModule_io_inputs_0),
    .io_inputs_1(regMaxVec_4_comparatorModule_io_inputs_1),
    .io_inputs_2(regMaxVec_4_comparatorModule_io_inputs_2),
    .io_inputs_3(regMaxVec_4_comparatorModule_io_inputs_3),
    .io_inputs_4(regMaxVec_4_comparatorModule_io_inputs_4),
    .io_result(regMaxVec_4_comparatorModule_io_result)
  );
  MultipleComparator_5 outResult_comparatorModule ( // @[multiple_comparator.scala 293:34]
    .clock(outResult_comparatorModule_clock),
    .io_start(outResult_comparatorModule_io_start),
    .io_inputs_0(outResult_comparatorModule_io_inputs_0),
    .io_inputs_1(outResult_comparatorModule_io_inputs_1),
    .io_inputs_2(outResult_comparatorModule_io_inputs_2),
    .io_inputs_3(outResult_comparatorModule_io_inputs_3),
    .io_inputs_4(outResult_comparatorModule_io_inputs_4),
    .io_result(outResult_comparatorModule_io_result)
  );
  assign io_outResultValid = 1'h0; // @[regular_fuzzification.scala 178:29 421:20]
  assign io_outResult = io_start ? outResult_result : 7'h0; // @[regular_fuzzification.scala 178:29 395:15 420:15]
  assign regMinVec_0_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_0_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_1_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_1_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_2_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_2_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_3_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_3_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_4_comparatorModule_io_in1 = regLutResultsVec_0; // @[comparator.scala 76:29]
  assign regMinVec_4_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_5_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_5_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_6_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_6_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_7_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_7_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_8_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_8_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_9_comparatorModule_io_in1 = regLutResultsVec_1; // @[comparator.scala 76:29]
  assign regMinVec_9_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_10_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_10_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_11_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_11_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_12_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_12_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_13_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_13_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_14_comparatorModule_io_in1 = regLutResultsVec_2; // @[comparator.scala 76:29]
  assign regMinVec_14_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_15_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_15_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_16_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_16_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_17_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_17_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_18_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_18_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_19_comparatorModule_io_in1 = regLutResultsVec_3; // @[comparator.scala 76:29]
  assign regMinVec_19_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMinVec_20_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_20_comparatorModule_io_in2 = regLutResultsVec_5; // @[comparator.scala 77:29]
  assign regMinVec_21_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_21_comparatorModule_io_in2 = regLutResultsVec_6; // @[comparator.scala 77:29]
  assign regMinVec_22_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_22_comparatorModule_io_in2 = regLutResultsVec_7; // @[comparator.scala 77:29]
  assign regMinVec_23_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_23_comparatorModule_io_in2 = regLutResultsVec_8; // @[comparator.scala 77:29]
  assign regMinVec_24_comparatorModule_io_in1 = regLutResultsVec_4; // @[comparator.scala 76:29]
  assign regMinVec_24_comparatorModule_io_in2 = regLutResultsVec_9; // @[comparator.scala 77:29]
  assign regMaxVec_0_comparatorModule_clock = clock;
  assign regMaxVec_0_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_0_comparatorModule_io_inputs_0 = regMinVec_0; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_0_comparatorModule_io_inputs_1 = regMinVec_1; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_0_comparatorModule_io_inputs_2 = regMinVec_2; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_0_comparatorModule_io_inputs_3 = regMinVec_5; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_1_comparatorModule_clock = clock;
  assign regMaxVec_1_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_1_comparatorModule_io_inputs_0 = regMinVec_3; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_1_comparatorModule_io_inputs_1 = regMinVec_4; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_1_comparatorModule_io_inputs_2 = regMinVec_6; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_1_comparatorModule_io_inputs_3 = regMinVec_7; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_1_comparatorModule_io_inputs_4 = regMinVec_8; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_1_comparatorModule_io_inputs_5 = regMinVec_10; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_2_comparatorModule_clock = clock;
  assign regMaxVec_2_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_2_comparatorModule_io_inputs_0 = regMinVec_9; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_2_comparatorModule_io_inputs_1 = regMinVec_11; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_2_comparatorModule_io_inputs_2 = regMinVec_12; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_2_comparatorModule_io_inputs_3 = regMinVec_15; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_3_comparatorModule_clock = clock;
  assign regMaxVec_3_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_3_comparatorModule_io_inputs_0 = regMinVec_13; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_3_comparatorModule_io_inputs_1 = regMinVec_14; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_3_comparatorModule_io_inputs_2 = regMinVec_16; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_3_comparatorModule_io_inputs_3 = regMinVec_17; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_3_comparatorModule_io_inputs_4 = regMinVec_20; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_3_comparatorModule_io_inputs_5 = regMinVec_21; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_4_comparatorModule_clock = clock;
  assign regMaxVec_4_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign regMaxVec_4_comparatorModule_io_inputs_0 = regMinVec_18; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_4_comparatorModule_io_inputs_1 = regMinVec_19; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_4_comparatorModule_io_inputs_2 = regMinVec_22; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_4_comparatorModule_io_inputs_3 = regMinVec_23; // @[regular_fuzzification.scala 323:15 326:30]
  assign regMaxVec_4_comparatorModule_io_inputs_4 = regMinVec_24; // @[regular_fuzzification.scala 323:15 326:30]
  assign outResult_comparatorModule_clock = clock;
  assign outResult_comparatorModule_io_start = io_start; // @[multiple_comparator.scala 309:31]
  assign outResult_comparatorModule_io_inputs_0 = regMaxVec_0; // @[regular_fuzzification.scala 378:11 385:40]
  assign outResult_comparatorModule_io_inputs_1 = regMaxVec_1; // @[regular_fuzzification.scala 378:11 385:40]
  assign outResult_comparatorModule_io_inputs_2 = regMaxVec_2; // @[regular_fuzzification.scala 378:11 385:40]
  assign outResult_comparatorModule_io_inputs_3 = regMaxVec_3; // @[regular_fuzzification.scala 378:11 385:40]
  assign outResult_comparatorModule_io_inputs_4 = regMaxVec_4; // @[regular_fuzzification.scala 378:11 385:40]
  always @(posedge clock) begin
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (10'h3ff == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_0 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fe == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_0 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fd == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_0 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_0 <= _GEN_1020;
      end
    end else begin
      regLutResultsVec_0 <= io_lutConnections_0; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (10'h3ff == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_1 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fe == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_1 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fd == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_1 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_1 <= _GEN_2044;
      end
    end else begin
      regLutResultsVec_1 <= io_lutConnections_1; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (10'h3ff == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_2 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fe == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_2 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fd == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_2 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_2 <= _GEN_3068;
      end
    end else begin
      regLutResultsVec_2 <= io_lutConnections_2; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (10'h3ff == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_3 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fe == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_3 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fd == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_3 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_3 <= _GEN_4092;
      end
    end else begin
      regLutResultsVec_3 <= io_lutConnections_3; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (10'h3ff == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_4 <= 7'h64; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fe == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_4 <= 7'h64; // @[regular_fuzzification.scala 194:38]
      end else if (10'h3fd == io_inputs_0) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_4 <= 7'h64; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_4 <= _GEN_5116;
      end
    end else begin
      regLutResultsVec_4 <= io_lutConnections_4; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (8'hff == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_5 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfe == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_5 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfd == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_5 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_5 <= _GEN_5372;
      end
    end else begin
      regLutResultsVec_5 <= io_lutConnections_5; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (8'hff == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_6 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfe == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_6 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfd == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_6 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_6 <= _GEN_5628;
      end
    end else begin
      regLutResultsVec_6 <= io_lutConnections_6; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (8'hff == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_7 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfe == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_7 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfd == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_7 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_7 <= _GEN_5884;
      end
    end else begin
      regLutResultsVec_7 <= io_lutConnections_7; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (8'hff == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_8 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfe == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_8 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfd == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_8 <= 7'h0; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_8 <= _GEN_6140;
      end
    end else begin
      regLutResultsVec_8 <= io_lutConnections_8; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (8'hff == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_9 <= 7'h64; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfe == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_9 <= 7'h64; // @[regular_fuzzification.scala 194:38]
      end else if (8'hfd == io_inputs_1[7:0]) begin // @[regular_fuzzification.scala 194:38]
        regLutResultsVec_9 <= 7'h64; // @[regular_fuzzification.scala 194:38]
      end else begin
        regLutResultsVec_9 <= _GEN_6396;
      end
    end else begin
      regLutResultsVec_9 <= io_lutConnections_9; // @[regular_fuzzification.scala 172:22]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_0_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_0 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_0 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_1_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_1 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_1 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_2_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_2 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_2 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_3_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_3 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_3 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_4_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_4 <= regLutResultsVec_0; // @[comparator.scala 101:14]
      end else begin
        regMinVec_4 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_5_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_5 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_5 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_6_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_6 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_6 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_7_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_7 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_7 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_8_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_8 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_8 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_9_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_9 <= regLutResultsVec_1; // @[comparator.scala 101:14]
      end else begin
        regMinVec_9 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_10_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_10 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_10 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_11_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_11 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_11 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_12_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_12 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_12 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_13_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_13 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_13 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_14_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_14 <= regLutResultsVec_2; // @[comparator.scala 101:14]
      end else begin
        regMinVec_14 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_15_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_15 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_15 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_16_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_16 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_16 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_17_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_17 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_17 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_18_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_18 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_18 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_19_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_19 <= regLutResultsVec_3; // @[comparator.scala 101:14]
      end else begin
        regMinVec_19 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_20_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_20 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_20 <= regLutResultsVec_5; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_21_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_21 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_21 <= regLutResultsVec_6; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_22_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_22 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_22 <= regLutResultsVec_7; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_23_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_23 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_23 <= regLutResultsVec_8; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      if (~regMinVec_24_maxMinOutput) begin // @[comparator.scala 100:40]
        regMinVec_24 <= regLutResultsVec_4; // @[comparator.scala 101:14]
      end else begin
        regMinVec_24 <= regLutResultsVec_9; // @[comparator.scala 103:14]
      end
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      regMaxVec_0 <= regMaxVec_0_result; // @[regular_fuzzification.scala 329:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      regMaxVec_1 <= regMaxVec_1_result; // @[regular_fuzzification.scala 329:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      regMaxVec_2 <= regMaxVec_2_result; // @[regular_fuzzification.scala 329:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      regMaxVec_3 <= regMaxVec_3_result; // @[regular_fuzzification.scala 329:39]
    end
    if (io_start) begin // @[regular_fuzzification.scala 178:29]
      regMaxVec_4 <= regMaxVec_4_result; // @[regular_fuzzification.scala 329:39]
    end
  end
endmodule
